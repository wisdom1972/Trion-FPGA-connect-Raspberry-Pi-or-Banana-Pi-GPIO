
//
// Verific Verilog Description of module top
//

module top (bscan_CAPTURE, bscan_DRCK, bscan_RESET, bscan_RUNTEST, bscan_SEL, 
            bscan_SHIFT, bscan_TCK, bscan_TDI, bscan_TMS, bscan_UPDATE, 
            bscan_TDO, clk, lock, raspi_gpiox8, freq_1sec_o, butten_o, 
            rasp0_i, rasp1_i, butten_i, led0_o, led1_o);
    input bscan_CAPTURE /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input bscan_DRCK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input bscan_RESET /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input bscan_RUNTEST /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input bscan_SEL /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input bscan_SHIFT /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input bscan_TCK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input bscan_TDI /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input bscan_TMS /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input bscan_UPDATE /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output bscan_TDO /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input clk /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input lock /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [7:0]raspi_gpiox8 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output freq_1sec_o /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output butten_o /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input rasp0_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input rasp1_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input butten_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output led0_o /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output led1_o /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    
    
    wire n24, n25, \cnt[0] , \edb_top/la0/la_run_trig , \edb_top/la0/la_trig_pattern[0] , 
        \edb_top/la0/la_run_trig_imdt , \edb_top/la0/la_stop_trig , \edb_top/la0/la_trig_mask[0] , 
        \edb_top/la0/address_counter[0] , n34, n35, n36, n37, \edb_top/la0/opcode[0] , 
        \edb_top/la0/bit_count[0] , n40, n41, \edb_top/la0/word_count[0] , 
        \edb_top/la0/data_out_shift_reg[0] , \edb_top/la0/module_state[0] , 
        \edb_top/la0/la_resetn_p1 , \edb_top/la0/cap_fifo_din[0] , \edb_top/la0/la_resetn , 
        \edb_top/la0/register_conn[64][0] , \edb_top/la0/register_conn[65][0] , 
        \edb_top/la0/register_conn[66][0] , \edb_top/la0/cap_fifo_din_p1[0] , 
        \edb_top/la0/cap_fifo_din_cu[0] , \edb_top/la0/cap_fifo_din_tu[0]_2 , 
        \edb_top/la0/internal_register_select[0] , \edb_top/la0/la_trig_pos[0] , 
        \edb_top/la0/la_trig_pattern[1] , \edb_top/la0/la_trig_mask[1] , 
        \edb_top/la0/la_trig_mask[2] , \edb_top/la0/la_trig_mask[3] , \edb_top/la0/la_trig_mask[4] , 
        \edb_top/la0/la_trig_mask[5] , \edb_top/la0/la_trig_mask[6] , \edb_top/la0/la_trig_mask[7] , 
        \edb_top/la0/la_trig_mask[8] , \edb_top/la0/la_trig_mask[9] , \edb_top/la0/la_trig_mask[10] , 
        \edb_top/la0/la_trig_mask[11] , \edb_top/la0/la_trig_mask[12] , 
        \edb_top/la0/la_trig_mask[13] , \edb_top/la0/la_trig_mask[14] , 
        \edb_top/la0/la_trig_mask[15] , \edb_top/la0/la_trig_mask[16] , 
        \edb_top/la0/la_trig_mask[17] , \edb_top/la0/la_trig_mask[18] , 
        \edb_top/la0/la_trig_mask[19] , \edb_top/la0/la_trig_mask[20] , 
        \edb_top/la0/la_trig_mask[21] , \edb_top/la0/la_trig_mask[22] , 
        \edb_top/la0/la_trig_mask[23] , \edb_top/la0/la_trig_mask[24] , 
        \edb_top/la0/la_trig_mask[25] , \edb_top/la0/la_trig_mask[26] , 
        \edb_top/la0/la_trig_mask[27] , \edb_top/la0/la_trig_mask[28] , 
        \edb_top/la0/la_trig_mask[29] , \edb_top/la0/la_trig_mask[30] , 
        \edb_top/la0/la_trig_mask[31] , \edb_top/la0/la_trig_mask[32] , 
        \edb_top/la0/la_trig_mask[33] , \edb_top/la0/la_trig_mask[34] , 
        \edb_top/la0/la_trig_mask[35] , \edb_top/la0/la_trig_mask[36] , 
        \edb_top/la0/la_trig_mask[37] , \edb_top/la0/la_trig_mask[38] , 
        \edb_top/la0/la_trig_mask[39] , \edb_top/la0/la_trig_mask[40] , 
        \edb_top/la0/la_trig_mask[41] , \edb_top/la0/la_trig_mask[42] , 
        \edb_top/la0/la_trig_mask[43] , \edb_top/la0/la_trig_mask[44] , 
        \edb_top/la0/la_trig_mask[45] , \edb_top/la0/la_trig_mask[46] , 
        \edb_top/la0/la_trig_mask[47] , \edb_top/la0/la_trig_mask[48] , 
        \edb_top/la0/la_trig_mask[49] , \edb_top/la0/la_trig_mask[50] , 
        \edb_top/la0/la_trig_mask[51] , \edb_top/la0/la_trig_mask[52] , 
        \edb_top/la0/la_trig_mask[53] , \edb_top/la0/la_trig_mask[54] , 
        \edb_top/la0/la_trig_mask[55] , \edb_top/la0/la_trig_mask[56] , 
        \edb_top/la0/la_trig_mask[57] , \edb_top/la0/la_trig_mask[58] , 
        \edb_top/la0/la_trig_mask[59] , \edb_top/la0/la_trig_mask[60] , 
        \edb_top/la0/la_trig_mask[61] , \edb_top/la0/la_trig_mask[62] , 
        \edb_top/la0/la_trig_mask[63] , \edb_top/la0/address_counter[1] , 
        \edb_top/la0/address_counter[2] , \edb_top/la0/address_counter[3] , 
        \edb_top/la0/address_counter[4] , \edb_top/la0/address_counter[5] , 
        \edb_top/la0/address_counter[6] , \edb_top/la0/address_counter[7] , 
        \edb_top/la0/address_counter[8] , \edb_top/la0/address_counter[9] , 
        \edb_top/la0/address_counter[10] , \edb_top/la0/address_counter[11] , 
        \edb_top/la0/address_counter[12] , \edb_top/la0/address_counter[13] , 
        \edb_top/la0/address_counter[14] , \edb_top/la0/address_counter[15] , 
        \edb_top/la0/address_counter[16] , \edb_top/la0/address_counter[17] , 
        \edb_top/la0/address_counter[18] , \edb_top/la0/address_counter[19] , 
        \edb_top/la0/address_counter[20] , \edb_top/la0/address_counter[21] , 
        \edb_top/la0/address_counter[22] , \edb_top/la0/address_counter[23] , 
        \edb_top/la0/address_counter[24] , \edb_top/la0/opcode[1] , \edb_top/la0/opcode[2] , 
        \edb_top/la0/opcode[3] , \edb_top/la0/bit_count[1] , \edb_top/la0/bit_count[2] , 
        \edb_top/la0/bit_count[3] , \edb_top/la0/bit_count[4] , \edb_top/la0/bit_count[5] , 
        \edb_top/la0/word_count[1] , \edb_top/la0/word_count[2] , \edb_top/la0/word_count[3] , 
        \edb_top/la0/word_count[4] , \edb_top/la0/word_count[5] , \edb_top/la0/word_count[6] , 
        \edb_top/la0/word_count[7] , \edb_top/la0/word_count[8] , \edb_top/la0/word_count[9] , 
        \edb_top/la0/word_count[10] , \edb_top/la0/word_count[11] , \edb_top/la0/word_count[12] , 
        \edb_top/la0/word_count[13] , \edb_top/la0/word_count[14] , \edb_top/la0/word_count[15] , 
        \edb_top/la0/data_out_shift_reg[1] , \edb_top/la0/data_out_shift_reg[2] , 
        \edb_top/la0/data_out_shift_reg[3] , \edb_top/la0/data_out_shift_reg[4] , 
        \edb_top/la0/data_out_shift_reg[5] , \edb_top/la0/data_out_shift_reg[6] , 
        \edb_top/la0/data_out_shift_reg[7] , \edb_top/la0/data_out_shift_reg[8] , 
        \edb_top/la0/data_out_shift_reg[9] , \edb_top/la0/data_out_shift_reg[10] , 
        \edb_top/la0/data_out_shift_reg[11] , \edb_top/la0/data_out_shift_reg[12] , 
        \edb_top/la0/data_out_shift_reg[13] , \edb_top/la0/data_out_shift_reg[14] , 
        \edb_top/la0/data_out_shift_reg[15] , \edb_top/la0/data_out_shift_reg[16] , 
        \edb_top/la0/data_out_shift_reg[17] , \edb_top/la0/data_out_shift_reg[18] , 
        \edb_top/la0/data_out_shift_reg[19] , \edb_top/la0/data_out_shift_reg[20] , 
        \edb_top/la0/data_out_shift_reg[21] , \edb_top/la0/data_out_shift_reg[22] , 
        \edb_top/la0/data_out_shift_reg[23] , \edb_top/la0/data_out_shift_reg[24] , 
        \edb_top/la0/data_out_shift_reg[25] , \edb_top/la0/data_out_shift_reg[26] , 
        \edb_top/la0/data_out_shift_reg[27] , \edb_top/la0/data_out_shift_reg[28] , 
        \edb_top/la0/data_out_shift_reg[29] , \edb_top/la0/data_out_shift_reg[30] , 
        \edb_top/la0/data_out_shift_reg[31] , \edb_top/la0/data_out_shift_reg[32] , 
        \edb_top/la0/data_out_shift_reg[33] , \edb_top/la0/data_out_shift_reg[34] , 
        \edb_top/la0/data_out_shift_reg[35] , \edb_top/la0/data_out_shift_reg[36] , 
        \edb_top/la0/data_out_shift_reg[37] , \edb_top/la0/data_out_shift_reg[38] , 
        \edb_top/la0/data_out_shift_reg[39] , \edb_top/la0/data_out_shift_reg[40] , 
        \edb_top/la0/data_out_shift_reg[41] , \edb_top/la0/data_out_shift_reg[42] , 
        \edb_top/la0/data_out_shift_reg[43] , \edb_top/la0/data_out_shift_reg[44] , 
        \edb_top/la0/data_out_shift_reg[45] , \edb_top/la0/data_out_shift_reg[46] , 
        \edb_top/la0/data_out_shift_reg[47] , \edb_top/la0/data_out_shift_reg[48] , 
        \edb_top/la0/data_out_shift_reg[49] , \edb_top/la0/data_out_shift_reg[50] , 
        \edb_top/la0/data_out_shift_reg[51] , \edb_top/la0/data_out_shift_reg[52] , 
        \edb_top/la0/data_out_shift_reg[53] , \edb_top/la0/data_out_shift_reg[54] , 
        \edb_top/la0/data_out_shift_reg[55] , \edb_top/la0/data_out_shift_reg[56] , 
        \edb_top/la0/data_out_shift_reg[57] , \edb_top/la0/data_out_shift_reg[58] , 
        \edb_top/la0/data_out_shift_reg[59] , \edb_top/la0/data_out_shift_reg[60] , 
        \edb_top/la0/data_out_shift_reg[61] , \edb_top/la0/data_out_shift_reg[62] , 
        \edb_top/la0/data_out_shift_reg[63] , \edb_top/la0/module_state[1] , 
        \edb_top/la0/module_state[2] , \edb_top/la0/module_state[3] , \edb_top/la0/crc_data_out[0] , 
        \edb_top/la0/crc_data_out[1] , \edb_top/la0/crc_data_out[2] , \edb_top/la0/crc_data_out[3] , 
        \edb_top/la0/crc_data_out[4] , \edb_top/la0/crc_data_out[5] , \edb_top/la0/crc_data_out[6] , 
        \edb_top/la0/crc_data_out[7] , \edb_top/la0/crc_data_out[8] , \edb_top/la0/crc_data_out[9] , 
        \edb_top/la0/crc_data_out[10] , \edb_top/la0/crc_data_out[11] , 
        \edb_top/la0/crc_data_out[12] , \edb_top/la0/crc_data_out[13] , 
        \edb_top/la0/crc_data_out[14] , \edb_top/la0/crc_data_out[15] , 
        \edb_top/la0/crc_data_out[16] , \edb_top/la0/crc_data_out[17] , 
        \edb_top/la0/crc_data_out[18] , \edb_top/la0/crc_data_out[19] , 
        \edb_top/la0/crc_data_out[20] , \edb_top/la0/crc_data_out[21] , 
        \edb_top/la0/crc_data_out[22] , \edb_top/la0/crc_data_out[23] , 
        \edb_top/la0/crc_data_out[24] , \edb_top/la0/crc_data_out[25] , 
        \edb_top/la0/crc_data_out[26] , \edb_top/la0/crc_data_out[27] , 
        \edb_top/la0/crc_data_out[28] , \edb_top/la0/crc_data_out[29] , 
        \edb_top/la0/crc_data_out[30] , \edb_top/la0/crc_data_out[31] , 
        \edb_top/la0/cap_fifo_din[1] , \edb_top/la0/cap_fifo_din[2] , \edb_top/la0/cap_fifo_din[3] , 
        \edb_top/la0/cap_fifo_din[4] , \edb_top/la0/cap_fifo_din[5] , \edb_top/la0/cap_fifo_din[6] , 
        \edb_top/la0/cap_fifo_din[7] , \edb_top/la0/register_conn[64][1] , 
        \edb_top/la0/register_conn[64][2] , \edb_top/la0/register_conn[65][1] , 
        \edb_top/la0/register_conn[65][2] , \edb_top/la0/register_conn[65][3] , 
        \edb_top/la0/register_conn[65][4] , \edb_top/la0/register_conn[65][5] , 
        \edb_top/la0/register_conn[65][6] , \edb_top/la0/register_conn[65][7] , 
        \edb_top/la0/register_conn[65][8] , \edb_top/la0/register_conn[65][9] , 
        \edb_top/la0/register_conn[65][10] , \edb_top/la0/register_conn[65][11] , 
        \edb_top/la0/register_conn[65][12] , \edb_top/la0/register_conn[65][13] , 
        \edb_top/la0/register_conn[65][14] , \edb_top/la0/register_conn[65][15] , 
        \edb_top/la0/register_conn[65][16] , \edb_top/la0/register_conn[65][17] , 
        \edb_top/la0/register_conn[65][18] , \edb_top/la0/register_conn[65][19] , 
        \edb_top/la0/register_conn[65][20] , \edb_top/la0/register_conn[65][21] , 
        \edb_top/la0/register_conn[65][22] , \edb_top/la0/register_conn[65][23] , 
        \edb_top/la0/register_conn[65][24] , \edb_top/la0/register_conn[65][25] , 
        \edb_top/la0/register_conn[65][26] , \edb_top/la0/register_conn[65][27] , 
        \edb_top/la0/register_conn[65][28] , \edb_top/la0/register_conn[65][29] , 
        \edb_top/la0/register_conn[65][30] , \edb_top/la0/register_conn[65][31] , 
        \edb_top/la0/register_conn[65][32] , \edb_top/la0/register_conn[65][33] , 
        \edb_top/la0/register_conn[65][34] , \edb_top/la0/register_conn[65][35] , 
        \edb_top/la0/register_conn[65][36] , \edb_top/la0/register_conn[65][37] , 
        \edb_top/la0/register_conn[65][38] , \edb_top/la0/register_conn[65][39] , 
        \edb_top/la0/register_conn[65][40] , \edb_top/la0/register_conn[65][41] , 
        \edb_top/la0/register_conn[65][42] , \edb_top/la0/register_conn[65][43] , 
        \edb_top/la0/register_conn[65][44] , \edb_top/la0/register_conn[65][45] , 
        \edb_top/la0/register_conn[65][46] , \edb_top/la0/register_conn[65][47] , 
        \edb_top/la0/register_conn[65][48] , \edb_top/la0/register_conn[65][49] , 
        \edb_top/la0/register_conn[65][50] , \edb_top/la0/register_conn[65][51] , 
        \edb_top/la0/register_conn[65][52] , \edb_top/la0/register_conn[65][53] , 
        \edb_top/la0/register_conn[65][54] , \edb_top/la0/register_conn[65][55] , 
        \edb_top/la0/register_conn[65][56] , \edb_top/la0/register_conn[65][57] , 
        \edb_top/la0/register_conn[65][58] , \edb_top/la0/register_conn[65][59] , 
        \edb_top/la0/register_conn[65][60] , \edb_top/la0/register_conn[65][61] , 
        \edb_top/la0/register_conn[65][62] , \edb_top/la0/register_conn[65][63] , 
        \edb_top/la0/register_conn[66][1] , \edb_top/la0/register_conn[66][2] , 
        \edb_top/la0/register_conn[66][3] , \edb_top/la0/register_conn[66][4] , 
        \edb_top/la0/register_conn[66][5] , \edb_top/la0/register_conn[66][6] , 
        \edb_top/la0/register_conn[66][7] , \edb_top/la0/register_conn[66][8] , 
        \edb_top/la0/register_conn[66][9] , \edb_top/la0/register_conn[66][10] , 
        \edb_top/la0/register_conn[66][11] , \edb_top/la0/register_conn[66][12] , 
        \edb_top/la0/register_conn[66][13] , \edb_top/la0/register_conn[66][14] , 
        \edb_top/la0/register_conn[66][15] , \edb_top/la0/register_conn[66][16] , 
        \edb_top/la0/register_conn[66][17] , \edb_top/la0/register_conn[66][18] , 
        \edb_top/la0/register_conn[66][19] , \edb_top/la0/register_conn[66][20] , 
        \edb_top/la0/register_conn[66][21] , \edb_top/la0/register_conn[66][22] , 
        \edb_top/la0/register_conn[66][23] , \edb_top/la0/register_conn[66][24] , 
        \edb_top/la0/register_conn[66][25] , \edb_top/la0/register_conn[66][26] , 
        \edb_top/la0/register_conn[66][27] , \edb_top/la0/register_conn[66][28] , 
        \edb_top/la0/register_conn[66][29] , \edb_top/la0/register_conn[66][30] , 
        \edb_top/la0/register_conn[66][31] , \edb_top/la0/register_conn[66][32] , 
        \edb_top/la0/register_conn[66][33] , \edb_top/la0/register_conn[66][34] , 
        \edb_top/la0/register_conn[66][35] , \edb_top/la0/register_conn[66][36] , 
        \edb_top/la0/register_conn[66][37] , \edb_top/la0/register_conn[66][38] , 
        \edb_top/la0/register_conn[66][39] , \edb_top/la0/register_conn[66][40] , 
        \edb_top/la0/register_conn[66][41] , \edb_top/la0/register_conn[66][42] , 
        \edb_top/la0/register_conn[66][43] , \edb_top/la0/register_conn[66][44] , 
        \edb_top/la0/register_conn[66][45] , \edb_top/la0/register_conn[66][46] , 
        \edb_top/la0/register_conn[66][47] , \edb_top/la0/register_conn[66][48] , 
        \edb_top/la0/register_conn[66][49] , \edb_top/la0/register_conn[66][50] , 
        \edb_top/la0/register_conn[66][51] , \edb_top/la0/register_conn[66][52] , 
        \edb_top/la0/register_conn[66][53] , \edb_top/la0/register_conn[66][54] , 
        \edb_top/la0/register_conn[66][55] , \edb_top/la0/register_conn[66][56] , 
        \edb_top/la0/register_conn[66][57] , \edb_top/la0/register_conn[66][58] , 
        \edb_top/la0/register_conn[66][59] , \edb_top/la0/register_conn[66][60] , 
        \edb_top/la0/register_conn[66][61] , \edb_top/la0/register_conn[66][62] , 
        \edb_top/la0/register_conn[66][63] , \edb_top/la0/cap_fifo_din_p1[1] , 
        \edb_top/la0/cap_fifo_din_p1[2] , \edb_top/la0/cap_fifo_din_p1[3] , 
        \edb_top/la0/cap_fifo_din_p1[4] , \edb_top/la0/cap_fifo_din_p1[5] , 
        \edb_top/la0/cap_fifo_din_p1[6] , \edb_top/la0/cap_fifo_din_p1[7] , 
        \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[0] , \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp3[0] , 
        \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp4[0] , \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp5[0] , 
        \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp6[0] , \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[0] , 
        \edb_top/la0/tu_data[0] , \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[1] , 
        \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[2] , \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[3] , 
        \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[4] , \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[5] , 
        \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[6] , \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[7] , 
        \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[1] , \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[2] , 
        \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[3] , \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[4] , 
        \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[5] , \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[6] , 
        \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[7] , \edb_top/la0/tu_trigger , 
        \edb_top/la0/cap_fifo_din_cu[1] , \edb_top/la0/cap_fifo_din_cu[2] , 
        \edb_top/la0/cap_fifo_din_cu[3] , \edb_top/la0/cap_fifo_din_cu[4] , 
        \edb_top/la0/cap_fifo_din_cu[5] , \edb_top/la0/cap_fifo_din_cu[6] , 
        \edb_top/la0/cap_fifo_din_cu[7] , \edb_top/la0/cap_fifo_din_tu[1]_2 , 
        \edb_top/la0/cap_fifo_din_tu[2]_2 , \edb_top/la0/cap_fifo_din_tu[3]_2 , 
        \edb_top/la0/cap_fifo_din_tu[4]_2 , \edb_top/la0/cap_fifo_din_tu[5]_2 , 
        \edb_top/la0/cap_fifo_din_tu[6]_2 , \edb_top/la0/cap_fifo_din_tu[7]_2 , 
        \edb_top/la0/la_biu_inst/run_trig_p2 , \edb_top/la0/la_biu_inst/run_trig_imdt_p1 , 
        \edb_top/la0/la_biu_inst/run_trig_imdt_p2 , \edb_top/la0/la_biu_inst/cap_buf_read_done_p1 , 
        \edb_top/la0/la_biu_inst/cap_buf_read_done_p2 , \edb_top/la0/la_biu_inst/cap_buf_read_done_p3 , 
        n456, n457, \edb_top/la0/la_biu_inst/pos_counter[12] , \edb_top/la0/register_conn[0][0] , 
        \edb_top/la0/la_biu_inst/pos_counter[2] , \edb_top/la0/la_biu_inst/pos_counter[1] , 
        \edb_top/la0/la_biu_inst/pos_counter[0] , \edb_top/la0/la_biu_inst/pos_counter[13] , 
        \edb_top/la0/la_biu_inst/pos_counter[16] , \edb_top/la0/la_biu_inst/pos_counter[11] , 
        \edb_top/la0/la_biu_inst/str_sync , \edb_top/la0/la_biu_inst/str_sync_wbff1 , 
        \edb_top/la0/la_biu_inst/pos_counter[15] , \edb_top/la0/la_biu_inst/pos_counter[10] , 
        \edb_top/la0/la_biu_inst/str_sync_wbff2 , \edb_top/la0/la_biu_inst/str_sync_wbff2q , 
        \edb_top/la0/la_biu_inst/rdy_sync , \edb_top/la0/la_biu_inst/pos_counter[14] , 
        \edb_top/la0/la_biu_inst/pos_counter[9] , \edb_top/la0/la_biu_inst/rdy_sync_tff1 , 
        \edb_top/la0/la_biu_inst/rdy_sync_tff2 , \edb_top/la0/la_biu_inst/rdy_sync_tff2q , 
        \edb_top/la0/la_biu_inst/pos_counter[8] , \edb_top/la0/la_biu_inst/pos_counter[7] , 
        \edb_top/la0/la_biu_inst/pos_counter[6] , \edb_top/la0/data_from_biu[0] , 
        \edb_top/la0/la_biu_inst/pos_counter[5] , \edb_top/la0/la_biu_inst/pos_counter[4] , 
        \edb_top/la0/la_biu_inst/axi_fsm_state[0] , \edb_top/la0/la_biu_inst/pos_counter[3] , 
        \edb_top/la0/la_biu_inst/run_trig_p1 , \edb_top/la0/biu_ready , 
        \edb_top/la0/register_conn[0][1] , \edb_top/la0/register_conn[0][2] , 
        \edb_top/la0/la_biu_inst/row_addr[0] , \edb_top/la0/la_biu_inst/row_addr[1] , 
        \edb_top/la0/la_biu_inst/row_addr[2] , \edb_top/la0/la_biu_inst/row_addr[3] , 
        \edb_top/la0/la_biu_inst/row_addr[4] , \edb_top/la0/la_biu_inst/row_addr[5] , 
        \edb_top/la0/la_biu_inst/row_addr[6] , \edb_top/la0/la_biu_inst/row_addr[7] , 
        \edb_top/la0/la_biu_inst/row_addr[8] , \edb_top/la0/la_biu_inst/row_addr[9] , 
        \edb_top/la0/data_from_biu[1] , \edb_top/la0/data_from_biu[2] , 
        \edb_top/la0/data_from_biu[3] , \edb_top/la0/data_from_biu[4] , 
        \edb_top/la0/data_from_biu[5] , \edb_top/la0/data_from_biu[6] , 
        \edb_top/la0/data_from_biu[7] , \edb_top/la0/la_biu_inst/axi_fsm_state[1] , 
        n508, n509, \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0] , 
        n511, n512, \edb_top/la0/la_biu_inst/swapped_data_out[0] , \edb_top/la0/la_biu_inst/swapped_data_out[1] , 
        \edb_top/la0/la_biu_inst/swapped_data_out[2] , \edb_top/la0/la_biu_inst/swapped_data_out[3] , 
        \edb_top/la0/la_biu_inst/swapped_data_out[4] , \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]_2 , 
        \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1] , \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2] , 
        \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3] , \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4] , 
        \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5] , \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6] , 
        \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7] , \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8] , 
        \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9] , \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10] , 
        \edb_top/la0/la_biu_inst/swapped_data_out[5] , \edb_top/la0/la_biu_inst/swapped_data_out[6] , 
        \edb_top/la0/la_biu_inst/swapped_data_out[7] , n532, n533, n534, 
        n535, \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]_2 , 
        \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]_2 , \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]_2 , 
        \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]_2 , \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]_2 , 
        \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]_2 , \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]_2 , 
        \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]_2 , \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]_2 , 
        \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , \edb_top/la0/internal_register_select[1] , 
        \edb_top/la0/internal_register_select[2] , \edb_top/la0/internal_register_select[3] , 
        \edb_top/la0/internal_register_select[4] , \edb_top/la0/internal_register_select[5] , 
        \edb_top/la0/internal_register_select[6] , \edb_top/la0/internal_register_select[7] , 
        \edb_top/la0/internal_register_select[8] , \edb_top/la0/internal_register_select[9] , 
        \edb_top/la0/internal_register_select[10] , \edb_top/la0/internal_register_select[11] , 
        \edb_top/la0/internal_register_select[12] , \edb_top/la0/la_trig_pos[1] , 
        \edb_top/la0/la_trig_pos[2] , \edb_top/la0/la_trig_pos[3] , \edb_top/la0/la_trig_pos[4] , 
        \edb_top/la0/la_trig_pos[5] , \edb_top/la0/la_trig_pos[6] , \edb_top/la0/la_trig_pos[7] , 
        \edb_top/la0/la_trig_pos[8] , \edb_top/la0/la_trig_pos[9] , \edb_top/la0/la_trig_pos[10] , 
        \edb_top/la0/la_trig_pos[11] , \edb_top/la0/la_trig_pos[12] , \edb_top/la0/la_trig_pos[13] , 
        \edb_top/la0/la_trig_pos[14] , \edb_top/la0/la_trig_pos[15] , \edb_top/la0/la_trig_pos[16] , 
        n574, n575, n576, n577, n578, n579, n580, n581, n582, 
        n583, n584, n585, n586, n587, n588, n589, n590, n591, 
        n592, n593, n594, n595, n596, n597, n598, n599, n600, 
        n601, n602, n603, n604, n605, n606, n607, n608, n609, 
        n610, n611, n612, n613, n614, n615, n616, n617, n618, 
        n619, n620, n621, n622, n623, n624, n625, n626, n627, 
        n628, n629, n630, n631, n632, n633, n634, n635, n636, 
        n637, n638, n639, n640, n641, n642, n643, n644, n645, 
        n646, n647, n648, n649, n650, n651, n652, n653, n654, 
        n655, n656, n657, n658, n659, n660, n661, n662, n663, 
        n664, n665, n666, n667, n668, n669, n670, n671, n672, 
        n673, n674, n675, n676, n677, n678, n679, n680, n681, 
        n682, n683, n684, n685, n686, n687, \edb_top/debug_hub_inst/module_id_reg[0] , 
        n689, \edb_top/edb_user_dr[0] , n691, n692, n693, n694, 
        n695, n696, n710, n712, n713, n714, n715, n716, n717, 
        n718, n719, n720, n721, n722, n723, n724, n725, n726, 
        n727, n728, n729, n730, n731, n732, n733, n734, n735, 
        n736, n737, n738, n739, n740, n741, n742, n743, n744, 
        n745, n746, n747, n748, n749, n750, n751, n752, n753, 
        n754, n755, n756, n757, n771, n773, n774, n775, n776, 
        n777, n778, n779, n780, n781, n782, n783, n784, n785, 
        n786, n787, n788, n789, n790, n791, n792, n793, n794, 
        n795, n796, n797, n798, n799, n800, n801, n802, n803, 
        n804, n805, n806, n807, n808, n809, n810, n811, n812, 
        n813, n814, n815, n816, n817, n818, n819, n820, n821, 
        n822, n823, n824, n825, n826, n827, n828, n829, n830, 
        n831, n832, n833, n834, n835, n836, n837, n838, n839, 
        \edb_top/debug_hub_inst/module_id_reg[1] , \edb_top/debug_hub_inst/module_id_reg[2] , 
        \edb_top/debug_hub_inst/module_id_reg[3] , n843, n844, n845, 
        n846, n847, n848, \edb_top/edb_user_dr[1] , \edb_top/edb_user_dr[2] , 
        \edb_top/edb_user_dr[3] , \edb_top/edb_user_dr[4] , \edb_top/edb_user_dr[5] , 
        \edb_top/edb_user_dr[6] , \edb_top/edb_user_dr[7] , \edb_top/edb_user_dr[8] , 
        \edb_top/edb_user_dr[9] , \edb_top/edb_user_dr[10] , \edb_top/edb_user_dr[11] , 
        \edb_top/edb_user_dr[12] , \edb_top/edb_user_dr[13] , \edb_top/edb_user_dr[14] , 
        \edb_top/edb_user_dr[15] , \edb_top/edb_user_dr[16] , \edb_top/edb_user_dr[17] , 
        \edb_top/edb_user_dr[18] , \edb_top/edb_user_dr[19] , \edb_top/edb_user_dr[20] , 
        \edb_top/edb_user_dr[21] , \edb_top/edb_user_dr[22] , \edb_top/edb_user_dr[23] , 
        \edb_top/edb_user_dr[24] , \edb_top/edb_user_dr[25] , \edb_top/edb_user_dr[26] , 
        \edb_top/edb_user_dr[27] , \edb_top/edb_user_dr[28] , \edb_top/edb_user_dr[29] , 
        \edb_top/edb_user_dr[30] , \edb_top/edb_user_dr[31] , \edb_top/edb_user_dr[32] , 
        \edb_top/edb_user_dr[33] , \edb_top/edb_user_dr[34] , \edb_top/edb_user_dr[35] , 
        \edb_top/edb_user_dr[36] , \edb_top/edb_user_dr[37] , \edb_top/edb_user_dr[38] , 
        \edb_top/edb_user_dr[39] , \edb_top/edb_user_dr[40] , \edb_top/edb_user_dr[41] , 
        \edb_top/edb_user_dr[42] , \edb_top/edb_user_dr[43] , \edb_top/edb_user_dr[44] , 
        \edb_top/edb_user_dr[45] , \edb_top/edb_user_dr[46] , \edb_top/edb_user_dr[47] , 
        \edb_top/edb_user_dr[48] , \edb_top/edb_user_dr[49] , \edb_top/edb_user_dr[50] , 
        \edb_top/edb_user_dr[51] , \edb_top/edb_user_dr[52] , \edb_top/edb_user_dr[53] , 
        \edb_top/edb_user_dr[54] , \edb_top/edb_user_dr[55] , \edb_top/edb_user_dr[56] , 
        \edb_top/edb_user_dr[57] , \edb_top/edb_user_dr[58] , \edb_top/edb_user_dr[59] , 
        \edb_top/edb_user_dr[60] , \edb_top/edb_user_dr[61] , \edb_top/edb_user_dr[62] , 
        \edb_top/edb_user_dr[63] , \edb_top/edb_user_dr[64] , \edb_top/edb_user_dr[65] , 
        \edb_top/edb_user_dr[66] , \edb_top/edb_user_dr[67] , \edb_top/edb_user_dr[68] , 
        \edb_top/edb_user_dr[69] , \edb_top/edb_user_dr[70] , \edb_top/edb_user_dr[71] , 
        \edb_top/edb_user_dr[72] , \edb_top/edb_user_dr[73] , \edb_top/edb_user_dr[74] , 
        \edb_top/edb_user_dr[75] , \edb_top/edb_user_dr[76] , \edb_top/edb_user_dr[77] , 
        \edb_top/edb_user_dr[78] , \edb_top/edb_user_dr[79] , \edb_top/edb_user_dr[80] , 
        \edb_top/edb_user_dr[81] , \cnt[1] , \cnt[2] , \cnt[3] , \cnt[4] , 
        \cnt[5] , \cnt[6] , \cnt[7] , \cnt[8] , \cnt[9] , \cnt[10] , 
        \cnt[11] , \cnt[12] , \cnt[13] , \cnt[14] , \cnt[15] , \cnt[16] , 
        \cnt[17] , \cnt[18] , \cnt[19] , \cnt[20] , \cnt[21] , \cnt[22] , 
        \cnt[23] , \cnt[24] , \cnt[25] , \cnt[26] , \cnt[27] , \cnt[28] , 
        \cnt[29] , \cnt[30] , n969, n972, n973, n975, n978, n979, 
        n980, n982, n983, n984, n986, n990, n991, n992, n994, 
        n995, n996, n997, n998, n1001, n1002, n1003, n1008, 
        n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, 
        n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, 
        n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, 
        n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, 
        n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, 
        n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, 
        n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, 
        n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, 
        n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, 
        n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, 
        n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, 
        n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, 
        n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, 
        n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, 
        n1193, n1194, n1195, n1196, n1197, n1199, n1200, n1201, 
        n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, 
        n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, 
        n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1239, 
        n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, 
        n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, 
        n1256, n1257, n1258, n1277, n1282, n1283, n1284, n1285, 
        n1286, n1287, n1288, n1289, n1290, n1292, n1293, n1294, 
        n1298, n1299, n1300, n1303, n1304, n1305, n1307, n1308, 
        n1309, n1310, n1311, n1313, n1314, n1315, n1331, n1335, 
        n1336, \edb_top/la0/la_biu_inst/fifo_with_read_inst/n136 , \edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] , 
        \edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , \edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
        \edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , \edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
        \edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , \edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
        \edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , \edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
        \edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , \edb_top/la0/la_biu_inst/fifo_with_read_inst/we , 
        n1514, n1517, \bscan_TCK~O , \clk_2~O , n2039, n2038, n1683, 
        n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, 
        n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, 
        n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, 
        n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, 
        n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, 
        n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, 
        n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, 
        n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, 
        n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, 
        n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, 
        n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, 
        n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, 
        n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, 
        n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, 
        n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, 
        n1804, n1805, n1806, n1807, n1815, n1816, n1817, n1818, 
        n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, 
        n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, 
        n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, 
        n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, 
        n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, 
        n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, 
        n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, 
        n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, 
        n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, 
        n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, 
        n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, 
        n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, 
        n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, 
        n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, 
        n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, 
        n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, 
        n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, 
        n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, 
        n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, 
        n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, 
        n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, 
        n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, 
        n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, 
        n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, 
        n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, 
        n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, 
        n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, 
        n2035, n2036, n2037;
    
    assign led0_o = rasp0_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    assign led1_o = rasp1_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    assign butten_o = butten_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    EFX_LUT4 LUT__2645 (.I0(n1683), .I1(bscan_CAPTURE), .O(n1684)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2645.LUTMASK = 16'h8888;
    EFX_FF \freq_1sec~FF  (.D(freq_1sec_o), .CE(n969), .CLK(\clk_2~O ), 
           .SR(lock), .Q(freq_1sec_o)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \freq_1sec~FF .CLK_POLARITY = 1'b1;
    defparam \freq_1sec~FF .CE_POLARITY = 1'b0;
    defparam \freq_1sec~FF .SR_POLARITY = 1'b0;
    defparam \freq_1sec~FF .D_POLARITY = 1'b0;
    defparam \freq_1sec~FF .SR_SYNC = 1'b1;
    defparam \freq_1sec~FF .SR_VALUE = 1'b0;
    defparam \freq_1sec~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \cnt[0]~FF  (.D(\cnt[0] ), .CE(1'b1), .CLK(\clk_2~O ), .SR(n972), 
           .Q(\cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \cnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \cnt[0]~FF .SR_POLARITY = 1'b1;
    defparam \cnt[0]~FF .D_POLARITY = 1'b0;
    defparam \cnt[0]~FF .SR_SYNC = 1'b1;
    defparam \cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_run_trig~FF  (.D(n973), .CE(n975), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/la_run_trig )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1073)
    defparam \edb_top/la0/la_run_trig~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_run_trig~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/la_run_trig~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_run_trig~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_run_trig~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_run_trig~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_run_trig~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_pattern[0]~FF  (.D(\edb_top/edb_user_dr[62] ), 
           .CE(n978), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_pattern[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1073)
    defparam \edb_top/la0/la_trig_pattern[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pattern[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pattern[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pattern[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pattern[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_pattern[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_pattern[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_run_trig_imdt~FF  (.D(n979), .CE(n975), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/la_run_trig_imdt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1073)
    defparam \edb_top/la0/la_run_trig_imdt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_run_trig_imdt~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/la_run_trig_imdt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_run_trig_imdt~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_run_trig_imdt~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_run_trig_imdt~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_run_trig_imdt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_stop_trig~FF  (.D(n980), .CE(n975), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/la_stop_trig )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1073)
    defparam \edb_top/la0/la_stop_trig~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_stop_trig~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/la_stop_trig~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_stop_trig~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_stop_trig~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_stop_trig~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_stop_trig~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[0]~FF  (.D(\edb_top/edb_user_dr[0] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/address_counter[0]~FF  (.D(n983), .CE(n984), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/address_counter[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1101)
    defparam \edb_top/la0/address_counter[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/address_counter[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/address_counter[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/opcode[0]~FF  (.D(\edb_top/edb_user_dr[77] ), .CE(n990), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/opcode[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1111)
    defparam \edb_top/la0/opcode[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/opcode[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/opcode[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/opcode[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/opcode[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/opcode[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/opcode[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/bit_count[0]~FF  (.D(n991), .CE(n992), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/bit_count[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1120)
    defparam \edb_top/la0/bit_count[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/bit_count[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/bit_count[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/bit_count[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/bit_count[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/bit_count[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/bit_count[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/word_count[0]~FF  (.D(n994), .CE(n995), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/word_count[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1138)
    defparam \edb_top/la0/word_count[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/word_count[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/word_count[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[0]~FF  (.D(n996), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/module_state[0]~FF  (.D(n998), .CE(1'b1), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/module_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1193)
    defparam \edb_top/la0/module_state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/module_state[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/module_state[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/module_state[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/module_state[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/module_state[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/module_state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_resetn_p1~FF  (.D(1'b1), .CE(1'b1), .CLK(\clk_2~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/la_resetn_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1504)
    defparam \edb_top/la0/la_resetn_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_resetn_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_resetn_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_resetn_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_resetn_p1~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_resetn_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_resetn_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/cap_fifo_din[0]~FF  (.D(butten_o), .CE(1'b1), .CLK(\clk_2~O ), 
           .SR(1'b0), .Q(\edb_top/la0/cap_fifo_din[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1526)
    defparam \edb_top/la0/cap_fifo_din[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/cap_fifo_din[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_resetn~FF  (.D(\edb_top/la0/la_resetn_p1 ), .CE(1'b1), 
           .CLK(\clk_2~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_resetn )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1504)
    defparam \edb_top/la0/la_resetn~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_resetn~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_resetn~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_resetn~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_resetn~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_resetn~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_resetn~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[64][0]~FF  (.D(\edb_top/edb_user_dr[0] ), 
           .CE(n1001), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[64][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1567)
    defparam \edb_top/la0/register_conn[64][0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[64][0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[64][0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[64][0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[64][0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[64][0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[64][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][0]~FF  (.D(\edb_top/edb_user_dr[0] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][0]~FF  (.D(\edb_top/edb_user_dr[0] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/cap_fifo_din_p1[0]~FF  (.D(\edb_top/la0/cap_fifo_din[0] ), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/cap_fifo_din_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1649)
    defparam \edb_top/la0/cap_fifo_din_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/cap_fifo_din_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/cap_fifo_din_cu[0]~FF  (.D(\edb_top/la0/cap_fifo_din_p1[0] ), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/cap_fifo_din_cu[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1649)
    defparam \edb_top/la0/cap_fifo_din_cu[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/cap_fifo_din_cu[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/cap_fifo_din_tu[0]~FF  (.D(\edb_top/la0/cap_fifo_din_cu[0] ), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/cap_fifo_din_tu[0]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1661)
    defparam \edb_top/la0/cap_fifo_din_tu[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/cap_fifo_din_tu[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/internal_register_select[0]~FF  (.D(\edb_top/edb_user_dr[64] ), 
           .CE(n1008), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/internal_register_select[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1036)
    defparam \edb_top/la0/internal_register_select[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/internal_register_select[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/internal_register_select[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_pos[0]~FF  (.D(\edb_top/edb_user_dr[45] ), 
           .CE(n978), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_pos[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1073)
    defparam \edb_top/la0/la_trig_pos[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_pos[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_pos[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_pattern[1]~FF  (.D(\edb_top/edb_user_dr[63] ), 
           .CE(n978), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_pattern[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1073)
    defparam \edb_top/la0/la_trig_pattern[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pattern[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pattern[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pattern[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pattern[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_pattern[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_pattern[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[1]~FF  (.D(\edb_top/edb_user_dr[1] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[2]~FF  (.D(\edb_top/edb_user_dr[2] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[3]~FF  (.D(\edb_top/edb_user_dr[3] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[4]~FF  (.D(\edb_top/edb_user_dr[4] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[5]~FF  (.D(\edb_top/edb_user_dr[5] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[6]~FF  (.D(\edb_top/edb_user_dr[6] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[7]~FF  (.D(\edb_top/edb_user_dr[7] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[8]~FF  (.D(\edb_top/edb_user_dr[8] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[9]~FF  (.D(\edb_top/edb_user_dr[9] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[10]~FF  (.D(\edb_top/edb_user_dr[10] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[11]~FF  (.D(\edb_top/edb_user_dr[11] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[12]~FF  (.D(\edb_top/edb_user_dr[12] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[13]~FF  (.D(\edb_top/edb_user_dr[13] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[14]~FF  (.D(\edb_top/edb_user_dr[14] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[15]~FF  (.D(\edb_top/edb_user_dr[15] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[16]~FF  (.D(\edb_top/edb_user_dr[16] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[17]~FF  (.D(\edb_top/edb_user_dr[17] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[18]~FF  (.D(\edb_top/edb_user_dr[18] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[19]~FF  (.D(\edb_top/edb_user_dr[19] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[20]~FF  (.D(\edb_top/edb_user_dr[20] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[21]~FF  (.D(\edb_top/edb_user_dr[21] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[22]~FF  (.D(\edb_top/edb_user_dr[22] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[23]~FF  (.D(\edb_top/edb_user_dr[23] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[24]~FF  (.D(\edb_top/edb_user_dr[24] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[25]~FF  (.D(\edb_top/edb_user_dr[25] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[26]~FF  (.D(\edb_top/edb_user_dr[26] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[27]~FF  (.D(\edb_top/edb_user_dr[27] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[28]~FF  (.D(\edb_top/edb_user_dr[28] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[29]~FF  (.D(\edb_top/edb_user_dr[29] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[30]~FF  (.D(\edb_top/edb_user_dr[30] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[31]~FF  (.D(\edb_top/edb_user_dr[31] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[32]~FF  (.D(\edb_top/edb_user_dr[32] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[32]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[33]~FF  (.D(\edb_top/edb_user_dr[33] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[33]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[34]~FF  (.D(\edb_top/edb_user_dr[34] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[34]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[35]~FF  (.D(\edb_top/edb_user_dr[35] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[35]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[36]~FF  (.D(\edb_top/edb_user_dr[36] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[36]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[37]~FF  (.D(\edb_top/edb_user_dr[37] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[37]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[38]~FF  (.D(\edb_top/edb_user_dr[38] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[38]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[38]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[39]~FF  (.D(\edb_top/edb_user_dr[39] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[39]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[39]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[40]~FF  (.D(\edb_top/edb_user_dr[40] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[40]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[41]~FF  (.D(\edb_top/edb_user_dr[41] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[41]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[42]~FF  (.D(\edb_top/edb_user_dr[42] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[42]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[43]~FF  (.D(\edb_top/edb_user_dr[43] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[43]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[43]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[44]~FF  (.D(\edb_top/edb_user_dr[44] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[44]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[44]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[45]~FF  (.D(\edb_top/edb_user_dr[45] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[45]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[45]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[46]~FF  (.D(\edb_top/edb_user_dr[46] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[46]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[46]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[47]~FF  (.D(\edb_top/edb_user_dr[47] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[47]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[47]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[48]~FF  (.D(\edb_top/edb_user_dr[48] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[48]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[48]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[49]~FF  (.D(\edb_top/edb_user_dr[49] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[49]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[49]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[50]~FF  (.D(\edb_top/edb_user_dr[50] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[50]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[50]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[51]~FF  (.D(\edb_top/edb_user_dr[51] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[51]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[51]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[52]~FF  (.D(\edb_top/edb_user_dr[52] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[52]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[52]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[53]~FF  (.D(\edb_top/edb_user_dr[53] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[53]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[53]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[54]~FF  (.D(\edb_top/edb_user_dr[54] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[54]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[54]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[55]~FF  (.D(\edb_top/edb_user_dr[55] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[55]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[55]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[56]~FF  (.D(\edb_top/edb_user_dr[56] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[56]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[56]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[57]~FF  (.D(\edb_top/edb_user_dr[57] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[57]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[57]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[58]~FF  (.D(\edb_top/edb_user_dr[58] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[58]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[58]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[59]~FF  (.D(\edb_top/edb_user_dr[59] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[59]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[59]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[60]~FF  (.D(\edb_top/edb_user_dr[60] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[60]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[60]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[61]~FF  (.D(\edb_top/edb_user_dr[61] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[61]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[61]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[62]~FF  (.D(\edb_top/edb_user_dr[62] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[62]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[62]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_mask[63]~FF  (.D(\edb_top/edb_user_dr[63] ), 
           .CE(n982), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_mask[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1083)
    defparam \edb_top/la0/la_trig_mask[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[63]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_mask[63]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_mask[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_mask[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/address_counter[1]~FF  (.D(n1071), .CE(n984), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/address_counter[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1101)
    defparam \edb_top/la0/address_counter[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/address_counter[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/address_counter[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/address_counter[2]~FF  (.D(n1072), .CE(n984), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/address_counter[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1101)
    defparam \edb_top/la0/address_counter[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/address_counter[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/address_counter[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/address_counter[3]~FF  (.D(n1073), .CE(n984), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/address_counter[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1101)
    defparam \edb_top/la0/address_counter[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/address_counter[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/address_counter[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/address_counter[4]~FF  (.D(n1074), .CE(n984), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/address_counter[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1101)
    defparam \edb_top/la0/address_counter[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/address_counter[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/address_counter[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/address_counter[5]~FF  (.D(n1075), .CE(n984), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/address_counter[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1101)
    defparam \edb_top/la0/address_counter[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/address_counter[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/address_counter[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/address_counter[6]~FF  (.D(n1076), .CE(n984), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/address_counter[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1101)
    defparam \edb_top/la0/address_counter[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/address_counter[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/address_counter[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/address_counter[7]~FF  (.D(n1077), .CE(n984), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/address_counter[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1101)
    defparam \edb_top/la0/address_counter[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/address_counter[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/address_counter[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/address_counter[8]~FF  (.D(n1078), .CE(n984), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/address_counter[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1101)
    defparam \edb_top/la0/address_counter[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/address_counter[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/address_counter[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/address_counter[9]~FF  (.D(n1079), .CE(n984), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/address_counter[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1101)
    defparam \edb_top/la0/address_counter[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/address_counter[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/address_counter[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/address_counter[10]~FF  (.D(n1080), .CE(n984), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/address_counter[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1101)
    defparam \edb_top/la0/address_counter[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/address_counter[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/address_counter[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/address_counter[11]~FF  (.D(n1081), .CE(n984), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/address_counter[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1101)
    defparam \edb_top/la0/address_counter[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/address_counter[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/address_counter[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/address_counter[12]~FF  (.D(n1082), .CE(n984), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/address_counter[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1101)
    defparam \edb_top/la0/address_counter[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/address_counter[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/address_counter[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/address_counter[13]~FF  (.D(n1083), .CE(n984), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/address_counter[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1101)
    defparam \edb_top/la0/address_counter[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/address_counter[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/address_counter[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/address_counter[14]~FF  (.D(n1084), .CE(n984), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/address_counter[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1101)
    defparam \edb_top/la0/address_counter[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/address_counter[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/address_counter[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/address_counter[15]~FF  (.D(n1085), .CE(n984), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/address_counter[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1101)
    defparam \edb_top/la0/address_counter[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/address_counter[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/address_counter[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/address_counter[16]~FF  (.D(n1086), .CE(n984), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/address_counter[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1101)
    defparam \edb_top/la0/address_counter[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/address_counter[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/address_counter[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/address_counter[17]~FF  (.D(n1087), .CE(n984), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/address_counter[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1101)
    defparam \edb_top/la0/address_counter[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/address_counter[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/address_counter[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/address_counter[18]~FF  (.D(n1088), .CE(n984), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/address_counter[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1101)
    defparam \edb_top/la0/address_counter[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/address_counter[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/address_counter[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/address_counter[19]~FF  (.D(n1089), .CE(n984), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/address_counter[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1101)
    defparam \edb_top/la0/address_counter[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/address_counter[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/address_counter[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/address_counter[20]~FF  (.D(n1090), .CE(n984), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/address_counter[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1101)
    defparam \edb_top/la0/address_counter[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/address_counter[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/address_counter[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/address_counter[21]~FF  (.D(n1091), .CE(n984), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/address_counter[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1101)
    defparam \edb_top/la0/address_counter[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/address_counter[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/address_counter[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/address_counter[22]~FF  (.D(n1092), .CE(n984), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/address_counter[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1101)
    defparam \edb_top/la0/address_counter[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/address_counter[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/address_counter[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/address_counter[23]~FF  (.D(n1093), .CE(n984), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/address_counter[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1101)
    defparam \edb_top/la0/address_counter[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/address_counter[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/address_counter[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/address_counter[24]~FF  (.D(n1094), .CE(n984), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/address_counter[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1101)
    defparam \edb_top/la0/address_counter[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/address_counter[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/address_counter[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/address_counter[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/opcode[1]~FF  (.D(\edb_top/edb_user_dr[78] ), .CE(n990), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/opcode[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1111)
    defparam \edb_top/la0/opcode[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/opcode[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/opcode[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/opcode[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/opcode[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/opcode[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/opcode[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/opcode[2]~FF  (.D(\edb_top/edb_user_dr[79] ), .CE(n990), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/opcode[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1111)
    defparam \edb_top/la0/opcode[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/opcode[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/opcode[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/opcode[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/opcode[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/opcode[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/opcode[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/opcode[3]~FF  (.D(\edb_top/edb_user_dr[80] ), .CE(n990), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/opcode[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1111)
    defparam \edb_top/la0/opcode[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/opcode[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/opcode[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/opcode[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/opcode[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/opcode[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/opcode[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/bit_count[1]~FF  (.D(n1105), .CE(n992), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/bit_count[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1120)
    defparam \edb_top/la0/bit_count[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/bit_count[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/bit_count[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/bit_count[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/bit_count[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/bit_count[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/bit_count[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/bit_count[2]~FF  (.D(n1106), .CE(n992), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/bit_count[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1120)
    defparam \edb_top/la0/bit_count[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/bit_count[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/bit_count[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/bit_count[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/bit_count[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/bit_count[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/bit_count[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/bit_count[3]~FF  (.D(n1107), .CE(n992), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/bit_count[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1120)
    defparam \edb_top/la0/bit_count[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/bit_count[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/bit_count[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/bit_count[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/bit_count[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/bit_count[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/bit_count[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/bit_count[4]~FF  (.D(n1108), .CE(n992), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/bit_count[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1120)
    defparam \edb_top/la0/bit_count[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/bit_count[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/bit_count[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/bit_count[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/bit_count[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/bit_count[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/bit_count[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/bit_count[5]~FF  (.D(n1109), .CE(n992), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/bit_count[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1120)
    defparam \edb_top/la0/bit_count[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/bit_count[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/bit_count[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/bit_count[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/bit_count[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/bit_count[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/bit_count[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/word_count[1]~FF  (.D(n1110), .CE(n995), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/word_count[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1138)
    defparam \edb_top/la0/word_count[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/word_count[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/word_count[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/word_count[2]~FF  (.D(n1111), .CE(n995), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/word_count[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1138)
    defparam \edb_top/la0/word_count[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/word_count[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/word_count[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/word_count[3]~FF  (.D(n1112), .CE(n995), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/word_count[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1138)
    defparam \edb_top/la0/word_count[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/word_count[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/word_count[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/word_count[4]~FF  (.D(n1113), .CE(n995), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/word_count[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1138)
    defparam \edb_top/la0/word_count[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/word_count[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/word_count[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/word_count[5]~FF  (.D(n1114), .CE(n995), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/word_count[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1138)
    defparam \edb_top/la0/word_count[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/word_count[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/word_count[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/word_count[6]~FF  (.D(n1115), .CE(n995), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/word_count[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1138)
    defparam \edb_top/la0/word_count[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/word_count[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/word_count[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/word_count[7]~FF  (.D(n1116), .CE(n995), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/word_count[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1138)
    defparam \edb_top/la0/word_count[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/word_count[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/word_count[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/word_count[8]~FF  (.D(n1117), .CE(n995), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/word_count[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1138)
    defparam \edb_top/la0/word_count[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/word_count[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/word_count[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/word_count[9]~FF  (.D(n1118), .CE(n995), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/word_count[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1138)
    defparam \edb_top/la0/word_count[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/word_count[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/word_count[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/word_count[10]~FF  (.D(n1119), .CE(n995), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/word_count[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1138)
    defparam \edb_top/la0/word_count[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/word_count[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/word_count[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/word_count[11]~FF  (.D(n1120), .CE(n995), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/word_count[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1138)
    defparam \edb_top/la0/word_count[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/word_count[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/word_count[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/word_count[12]~FF  (.D(n1121), .CE(n995), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/word_count[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1138)
    defparam \edb_top/la0/word_count[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/word_count[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/word_count[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/word_count[13]~FF  (.D(n1122), .CE(n995), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/word_count[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1138)
    defparam \edb_top/la0/word_count[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/word_count[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/word_count[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/word_count[14]~FF  (.D(n1123), .CE(n995), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/word_count[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1138)
    defparam \edb_top/la0/word_count[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/word_count[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/word_count[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/word_count[15]~FF  (.D(n1124), .CE(n995), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/word_count[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1138)
    defparam \edb_top/la0/word_count[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/word_count[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/word_count[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/word_count[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[1]~FF  (.D(n1125), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[2]~FF  (.D(n1126), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[3]~FF  (.D(n1127), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[4]~FF  (.D(n1128), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[5]~FF  (.D(n1129), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[6]~FF  (.D(n1130), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[7]~FF  (.D(n1131), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[8]~FF  (.D(n1132), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[9]~FF  (.D(n1133), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[10]~FF  (.D(n1134), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[11]~FF  (.D(n1135), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[11]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[12]~FF  (.D(n1136), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[12]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[13]~FF  (.D(n1137), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[13]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[14]~FF  (.D(n1138), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[14]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[15]~FF  (.D(n1139), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[15]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[16]~FF  (.D(n1140), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[16]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[17]~FF  (.D(n1141), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[17]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[18]~FF  (.D(n1142), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[18]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[19]~FF  (.D(n1143), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[19]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[20]~FF  (.D(n1144), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[20]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[21]~FF  (.D(n1145), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[21]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[22]~FF  (.D(n1146), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[22]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[23]~FF  (.D(n1147), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[23]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[24]~FF  (.D(n1148), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[24]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[25]~FF  (.D(n1149), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[25]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[26]~FF  (.D(n1150), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[26]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[27]~FF  (.D(n1151), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[27]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[28]~FF  (.D(n1152), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[28]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[29]~FF  (.D(n1153), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[29]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[30]~FF  (.D(n1154), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[30]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[31]~FF  (.D(n1155), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[31]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[32]~FF  (.D(n1156), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[32]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[32]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[33]~FF  (.D(n1157), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[33]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[33]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[34]~FF  (.D(n1158), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[34]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[34]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[35]~FF  (.D(n1159), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[35]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[35]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[36]~FF  (.D(n1160), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[36]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[36]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[37]~FF  (.D(n1161), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[37]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[37]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[38]~FF  (.D(n1162), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[38]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[38]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[39]~FF  (.D(n1163), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[39]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[39]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[40]~FF  (.D(n1164), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[40]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[40]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[41]~FF  (.D(n1165), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[41]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[41]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[42]~FF  (.D(n1166), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[42]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[42]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[43]~FF  (.D(n1167), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[43]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[43]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[44]~FF  (.D(n1168), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[44]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[44]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[45]~FF  (.D(n1169), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[45]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[45]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[46]~FF  (.D(n1170), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[46]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[46]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[47]~FF  (.D(n1171), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[47]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[47]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[48]~FF  (.D(n1172), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[48]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[48]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[49]~FF  (.D(n1173), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[49]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[49]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[50]~FF  (.D(n1174), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[50]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[50]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[51]~FF  (.D(n1175), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[51]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[51]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[52]~FF  (.D(n1176), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[52]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[52]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[53]~FF  (.D(n1177), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[53]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[53]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[54]~FF  (.D(n1178), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[54]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[54]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[55]~FF  (.D(n1179), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[55]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[55]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[56]~FF  (.D(n1180), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[56]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[56]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[57]~FF  (.D(n1181), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[57]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[57]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[58]~FF  (.D(n1182), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[58]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[58]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[59]~FF  (.D(n1183), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[59]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[59]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[60]~FF  (.D(n1184), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[60]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[60]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[61]~FF  (.D(n1185), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[61]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[61]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[62]~FF  (.D(n1186), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[62]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[62]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/data_out_shift_reg[63]~FF  (.D(n1187), .CE(n997), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/data_out_shift_reg[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1151)
    defparam \edb_top/la0/data_out_shift_reg[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[63]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/data_out_shift_reg[63]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/data_out_shift_reg[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/module_state[1]~FF  (.D(n1188), .CE(1'b1), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/module_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1193)
    defparam \edb_top/la0/module_state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/module_state[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/module_state[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/module_state[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/module_state[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/module_state[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/module_state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/module_state[2]~FF  (.D(n1189), .CE(1'b1), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/module_state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1193)
    defparam \edb_top/la0/module_state[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/module_state[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/module_state[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/module_state[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/module_state[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/module_state[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/module_state[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/module_state[3]~FF  (.D(n1190), .CE(1'b1), .CLK(\bscan_TCK~O ), 
           .SR(bscan_RESET), .Q(\edb_top/la0/module_state[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1193)
    defparam \edb_top/la0/module_state[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/module_state[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/module_state[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/module_state[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/module_state[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/module_state[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/module_state[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[0]~FF  (.D(n1191), 
           .CE(n1192), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/crc_data_out[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(234)
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[0]~FF .SR_VALUE = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[1]~FF  (.D(n1193), 
           .CE(n1192), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/crc_data_out[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(234)
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[1]~FF .SR_VALUE = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[2]~FF  (.D(n1194), 
           .CE(n1192), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/crc_data_out[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(234)
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[2]~FF .SR_VALUE = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[3]~FF  (.D(n1195), 
           .CE(n1192), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/crc_data_out[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(234)
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[3]~FF .SR_VALUE = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[4]~FF  (.D(n1196), 
           .CE(n1192), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/crc_data_out[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(234)
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[4]~FF .SR_VALUE = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[5]~FF  (.D(n1197), 
           .CE(n1192), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/crc_data_out[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(234)
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[5]~FF .SR_VALUE = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[6]~FF  (.D(n1199), 
           .CE(n1192), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/crc_data_out[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(234)
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[6]~FF .SR_VALUE = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[7]~FF  (.D(n1200), 
           .CE(n1192), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/crc_data_out[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(234)
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[7]~FF .SR_VALUE = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[8]~FF  (.D(n1201), 
           .CE(n1192), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/crc_data_out[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(234)
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[8]~FF .SR_VALUE = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[9]~FF  (.D(n1202), 
           .CE(n1192), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/crc_data_out[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(234)
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[9]~FF .SR_VALUE = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[10]~FF  (.D(n1203), 
           .CE(n1192), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/crc_data_out[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(234)
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[10]~FF .SR_VALUE = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[11]~FF  (.D(n1204), 
           .CE(n1192), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/crc_data_out[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(234)
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[11]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[11]~FF .SR_VALUE = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[12]~FF  (.D(n1205), 
           .CE(n1192), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/crc_data_out[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(234)
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[12]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[12]~FF .SR_VALUE = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[13]~FF  (.D(n1206), 
           .CE(n1192), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/crc_data_out[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(234)
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[13]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[13]~FF .SR_VALUE = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[14]~FF  (.D(n1207), 
           .CE(n1192), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/crc_data_out[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(234)
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[14]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[14]~FF .SR_VALUE = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[15]~FF  (.D(n1208), 
           .CE(n1192), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/crc_data_out[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(234)
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[15]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[15]~FF .SR_VALUE = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[16]~FF  (.D(n1209), 
           .CE(n1192), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/crc_data_out[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(234)
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[16]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[16]~FF .SR_VALUE = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[17]~FF  (.D(n1210), 
           .CE(n1192), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/crc_data_out[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(234)
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[17]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[17]~FF .SR_VALUE = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[18]~FF  (.D(n1211), 
           .CE(n1192), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/crc_data_out[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(234)
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[18]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[18]~FF .SR_VALUE = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[19]~FF  (.D(n1212), 
           .CE(n1192), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/crc_data_out[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(234)
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[19]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[19]~FF .SR_VALUE = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[20]~FF  (.D(n1213), 
           .CE(n1192), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/crc_data_out[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(234)
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[20]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[20]~FF .SR_VALUE = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[21]~FF  (.D(n1214), 
           .CE(n1192), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/crc_data_out[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(234)
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[21]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[21]~FF .SR_VALUE = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[22]~FF  (.D(n1215), 
           .CE(n1192), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/crc_data_out[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(234)
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[22]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[22]~FF .SR_VALUE = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[23]~FF  (.D(n1216), 
           .CE(n1192), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/crc_data_out[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(234)
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[23]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[23]~FF .SR_VALUE = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[24]~FF  (.D(n1217), 
           .CE(n1192), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/crc_data_out[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(234)
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[24]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[24]~FF .SR_VALUE = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[25]~FF  (.D(n1218), 
           .CE(n1192), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/crc_data_out[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(234)
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[25]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[25]~FF .SR_VALUE = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[26]~FF  (.D(n1219), 
           .CE(n1192), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/crc_data_out[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(234)
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[26]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[26]~FF .SR_VALUE = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[27]~FF  (.D(n1220), 
           .CE(n1192), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/crc_data_out[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(234)
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[27]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[27]~FF .SR_VALUE = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[28]~FF  (.D(n1221), 
           .CE(n1192), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/crc_data_out[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(234)
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[28]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[28]~FF .SR_VALUE = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[29]~FF  (.D(n1222), 
           .CE(n1192), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/crc_data_out[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(234)
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[29]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[29]~FF .SR_VALUE = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[30]~FF  (.D(n1223), 
           .CE(n1192), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/crc_data_out[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(234)
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[30]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[30]~FF .SR_VALUE = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[31]~FF  (.D(n1224), 
           .CE(n1192), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/crc_data_out[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(234)
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[31]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[31]~FF .SR_VALUE = 1'b1;
    defparam \edb_top/la0/axi_crc_i/edb_top/la0/crc_data_out[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/cap_fifo_din[1]~FF  (.D(raspi_gpiox8[0]), .CE(1'b1), 
           .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/cap_fifo_din[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1526)
    defparam \edb_top/la0/cap_fifo_din[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/cap_fifo_din[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/cap_fifo_din[2]~FF  (.D(raspi_gpiox8[1]), .CE(1'b1), 
           .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/cap_fifo_din[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1526)
    defparam \edb_top/la0/cap_fifo_din[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/cap_fifo_din[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/cap_fifo_din[3]~FF  (.D(raspi_gpiox8[2]), .CE(1'b1), 
           .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/cap_fifo_din[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1526)
    defparam \edb_top/la0/cap_fifo_din[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/cap_fifo_din[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/cap_fifo_din[4]~FF  (.D(raspi_gpiox8[3]), .CE(1'b1), 
           .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/cap_fifo_din[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1526)
    defparam \edb_top/la0/cap_fifo_din[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/cap_fifo_din[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/cap_fifo_din[5]~FF  (.D(raspi_gpiox8[4]), .CE(1'b1), 
           .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/cap_fifo_din[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1526)
    defparam \edb_top/la0/cap_fifo_din[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/cap_fifo_din[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/cap_fifo_din[6]~FF  (.D(raspi_gpiox8[5]), .CE(1'b1), 
           .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/cap_fifo_din[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1526)
    defparam \edb_top/la0/cap_fifo_din[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/cap_fifo_din[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/cap_fifo_din[7]~FF  (.D(raspi_gpiox8[6]), .CE(1'b1), 
           .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/cap_fifo_din[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1526)
    defparam \edb_top/la0/cap_fifo_din[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/cap_fifo_din[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/cap_fifo_din[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[64][1]~FF  (.D(\edb_top/edb_user_dr[1] ), 
           .CE(n1001), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[64][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1567)
    defparam \edb_top/la0/register_conn[64][1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[64][1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[64][1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[64][1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[64][1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[64][1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[64][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[64][2]~FF  (.D(\edb_top/edb_user_dr[2] ), 
           .CE(n1001), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[64][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1567)
    defparam \edb_top/la0/register_conn[64][2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[64][2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[64][2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[64][2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[64][2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[64][2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[64][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][1]~FF  (.D(\edb_top/edb_user_dr[1] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][2]~FF  (.D(\edb_top/edb_user_dr[2] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][3]~FF  (.D(\edb_top/edb_user_dr[3] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][4]~FF  (.D(\edb_top/edb_user_dr[4] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][5]~FF  (.D(\edb_top/edb_user_dr[5] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][6]~FF  (.D(\edb_top/edb_user_dr[6] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][7]~FF  (.D(\edb_top/edb_user_dr[7] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][8]~FF  (.D(\edb_top/edb_user_dr[8] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][9]~FF  (.D(\edb_top/edb_user_dr[9] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][10]~FF  (.D(\edb_top/edb_user_dr[10] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][11]~FF  (.D(\edb_top/edb_user_dr[11] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][12]~FF  (.D(\edb_top/edb_user_dr[12] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][13]~FF  (.D(\edb_top/edb_user_dr[13] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][14]~FF  (.D(\edb_top/edb_user_dr[14] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][15]~FF  (.D(\edb_top/edb_user_dr[15] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][16]~FF  (.D(\edb_top/edb_user_dr[16] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][17]~FF  (.D(\edb_top/edb_user_dr[17] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][18]~FF  (.D(\edb_top/edb_user_dr[18] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][19]~FF  (.D(\edb_top/edb_user_dr[19] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][20]~FF  (.D(\edb_top/edb_user_dr[20] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][21]~FF  (.D(\edb_top/edb_user_dr[21] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][22]~FF  (.D(\edb_top/edb_user_dr[22] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][23]~FF  (.D(\edb_top/edb_user_dr[23] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][24]~FF  (.D(\edb_top/edb_user_dr[24] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][25]~FF  (.D(\edb_top/edb_user_dr[25] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][26]~FF  (.D(\edb_top/edb_user_dr[26] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][27]~FF  (.D(\edb_top/edb_user_dr[27] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][28]~FF  (.D(\edb_top/edb_user_dr[28] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][29]~FF  (.D(\edb_top/edb_user_dr[29] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][30]~FF  (.D(\edb_top/edb_user_dr[30] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][31]~FF  (.D(\edb_top/edb_user_dr[31] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][32]~FF  (.D(\edb_top/edb_user_dr[32] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][32]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][33]~FF  (.D(\edb_top/edb_user_dr[33] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][33]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][34]~FF  (.D(\edb_top/edb_user_dr[34] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][34]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][35]~FF  (.D(\edb_top/edb_user_dr[35] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][35]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][36]~FF  (.D(\edb_top/edb_user_dr[36] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][36]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][37]~FF  (.D(\edb_top/edb_user_dr[37] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][37]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][38]~FF  (.D(\edb_top/edb_user_dr[38] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][38]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][38]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][39]~FF  (.D(\edb_top/edb_user_dr[39] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][39]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][39]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][40]~FF  (.D(\edb_top/edb_user_dr[40] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][40]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][41]~FF  (.D(\edb_top/edb_user_dr[41] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][41]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][42]~FF  (.D(\edb_top/edb_user_dr[42] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][42]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][43]~FF  (.D(\edb_top/edb_user_dr[43] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][43]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][43]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][44]~FF  (.D(\edb_top/edb_user_dr[44] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][44]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][44]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][45]~FF  (.D(\edb_top/edb_user_dr[45] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][45]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][45]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][46]~FF  (.D(\edb_top/edb_user_dr[46] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][46]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][46]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][47]~FF  (.D(\edb_top/edb_user_dr[47] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][47]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][47]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][48]~FF  (.D(\edb_top/edb_user_dr[48] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][48]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][48]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][49]~FF  (.D(\edb_top/edb_user_dr[49] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][49]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][49]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][50]~FF  (.D(\edb_top/edb_user_dr[50] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][50]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][50]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][51]~FF  (.D(\edb_top/edb_user_dr[51] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][51]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][51]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][52]~FF  (.D(\edb_top/edb_user_dr[52] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][52]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][52]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][53]~FF  (.D(\edb_top/edb_user_dr[53] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][53]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][53]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][54]~FF  (.D(\edb_top/edb_user_dr[54] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][54]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][54]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][55]~FF  (.D(\edb_top/edb_user_dr[55] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][55]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][55]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][56]~FF  (.D(\edb_top/edb_user_dr[56] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][56]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][56]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][57]~FF  (.D(\edb_top/edb_user_dr[57] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][57]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][57]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][58]~FF  (.D(\edb_top/edb_user_dr[58] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][58]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][58]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][59]~FF  (.D(\edb_top/edb_user_dr[59] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][59]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][59]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][60]~FF  (.D(\edb_top/edb_user_dr[60] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][60]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][60]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][61]~FF  (.D(\edb_top/edb_user_dr[61] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][61]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][61]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][62]~FF  (.D(\edb_top/edb_user_dr[62] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][62]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][62]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[65][63]~FF  (.D(\edb_top/edb_user_dr[63] ), 
           .CE(n1002), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[65][63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[65][63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][63]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[65][63]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[65][63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[65][63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][1]~FF  (.D(\edb_top/edb_user_dr[1] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][2]~FF  (.D(\edb_top/edb_user_dr[2] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][3]~FF  (.D(\edb_top/edb_user_dr[3] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][4]~FF  (.D(\edb_top/edb_user_dr[4] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][5]~FF  (.D(\edb_top/edb_user_dr[5] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][6]~FF  (.D(\edb_top/edb_user_dr[6] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][7]~FF  (.D(\edb_top/edb_user_dr[7] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][8]~FF  (.D(\edb_top/edb_user_dr[8] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][9]~FF  (.D(\edb_top/edb_user_dr[9] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][10]~FF  (.D(\edb_top/edb_user_dr[10] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][11]~FF  (.D(\edb_top/edb_user_dr[11] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][12]~FF  (.D(\edb_top/edb_user_dr[12] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][13]~FF  (.D(\edb_top/edb_user_dr[13] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][14]~FF  (.D(\edb_top/edb_user_dr[14] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][15]~FF  (.D(\edb_top/edb_user_dr[15] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][16]~FF  (.D(\edb_top/edb_user_dr[16] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][17]~FF  (.D(\edb_top/edb_user_dr[17] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][18]~FF  (.D(\edb_top/edb_user_dr[18] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][19]~FF  (.D(\edb_top/edb_user_dr[19] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][20]~FF  (.D(\edb_top/edb_user_dr[20] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][21]~FF  (.D(\edb_top/edb_user_dr[21] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][22]~FF  (.D(\edb_top/edb_user_dr[22] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][23]~FF  (.D(\edb_top/edb_user_dr[23] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][24]~FF  (.D(\edb_top/edb_user_dr[24] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][25]~FF  (.D(\edb_top/edb_user_dr[25] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][26]~FF  (.D(\edb_top/edb_user_dr[26] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][27]~FF  (.D(\edb_top/edb_user_dr[27] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][28]~FF  (.D(\edb_top/edb_user_dr[28] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][29]~FF  (.D(\edb_top/edb_user_dr[29] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][30]~FF  (.D(\edb_top/edb_user_dr[30] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][31]~FF  (.D(\edb_top/edb_user_dr[31] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][32]~FF  (.D(\edb_top/edb_user_dr[32] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][32]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][33]~FF  (.D(\edb_top/edb_user_dr[33] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][33]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][34]~FF  (.D(\edb_top/edb_user_dr[34] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][34]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][35]~FF  (.D(\edb_top/edb_user_dr[35] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][35]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][36]~FF  (.D(\edb_top/edb_user_dr[36] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][36]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][37]~FF  (.D(\edb_top/edb_user_dr[37] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][37]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][38]~FF  (.D(\edb_top/edb_user_dr[38] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][38]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][38]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][39]~FF  (.D(\edb_top/edb_user_dr[39] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][39]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][39]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][40]~FF  (.D(\edb_top/edb_user_dr[40] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][40]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][41]~FF  (.D(\edb_top/edb_user_dr[41] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][41]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][42]~FF  (.D(\edb_top/edb_user_dr[42] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][42]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][43]~FF  (.D(\edb_top/edb_user_dr[43] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][43]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][43]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][44]~FF  (.D(\edb_top/edb_user_dr[44] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][44]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][44]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][45]~FF  (.D(\edb_top/edb_user_dr[45] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][45]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][45]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][46]~FF  (.D(\edb_top/edb_user_dr[46] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][46]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][46]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][47]~FF  (.D(\edb_top/edb_user_dr[47] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][47]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][47]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][48]~FF  (.D(\edb_top/edb_user_dr[48] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][48]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][48]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][49]~FF  (.D(\edb_top/edb_user_dr[49] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][49]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][49]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][50]~FF  (.D(\edb_top/edb_user_dr[50] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][50]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][50]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][51]~FF  (.D(\edb_top/edb_user_dr[51] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][51]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][51]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][52]~FF  (.D(\edb_top/edb_user_dr[52] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][52]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][52]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][53]~FF  (.D(\edb_top/edb_user_dr[53] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][53]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][53]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][54]~FF  (.D(\edb_top/edb_user_dr[54] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][54]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][54]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][55]~FF  (.D(\edb_top/edb_user_dr[55] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][55]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][55]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][56]~FF  (.D(\edb_top/edb_user_dr[56] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][56]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][56]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][57]~FF  (.D(\edb_top/edb_user_dr[57] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][57]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][57]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][58]~FF  (.D(\edb_top/edb_user_dr[58] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][58]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][58]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][59]~FF  (.D(\edb_top/edb_user_dr[59] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][59]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][59]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][60]~FF  (.D(\edb_top/edb_user_dr[60] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][60]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][60]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][61]~FF  (.D(\edb_top/edb_user_dr[61] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][61]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][61]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][62]~FF  (.D(\edb_top/edb_user_dr[62] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][62]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][62]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/register_conn[66][63]~FF  (.D(\edb_top/edb_user_dr[63] ), 
           .CE(n1003), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/register_conn[66][63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1582)
    defparam \edb_top/la0/register_conn[66][63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][63]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/register_conn[66][63]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/register_conn[66][63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/register_conn[66][63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/cap_fifo_din_p1[1]~FF  (.D(\edb_top/la0/cap_fifo_din[1] ), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/cap_fifo_din_p1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1649)
    defparam \edb_top/la0/cap_fifo_din_p1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/cap_fifo_din_p1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/cap_fifo_din_p1[2]~FF  (.D(\edb_top/la0/cap_fifo_din[2] ), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/cap_fifo_din_p1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1649)
    defparam \edb_top/la0/cap_fifo_din_p1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/cap_fifo_din_p1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/cap_fifo_din_p1[3]~FF  (.D(\edb_top/la0/cap_fifo_din[3] ), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/cap_fifo_din_p1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1649)
    defparam \edb_top/la0/cap_fifo_din_p1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/cap_fifo_din_p1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/cap_fifo_din_p1[4]~FF  (.D(\edb_top/la0/cap_fifo_din[4] ), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/cap_fifo_din_p1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1649)
    defparam \edb_top/la0/cap_fifo_din_p1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/cap_fifo_din_p1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/cap_fifo_din_p1[5]~FF  (.D(\edb_top/la0/cap_fifo_din[5] ), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/cap_fifo_din_p1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1649)
    defparam \edb_top/la0/cap_fifo_din_p1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/cap_fifo_din_p1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/cap_fifo_din_p1[6]~FF  (.D(\edb_top/la0/cap_fifo_din[6] ), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/cap_fifo_din_p1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1649)
    defparam \edb_top/la0/cap_fifo_din_p1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/cap_fifo_din_p1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/cap_fifo_din_p1[7]~FF  (.D(\edb_top/la0/cap_fifo_din[7] ), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/cap_fifo_din_p1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1649)
    defparam \edb_top/la0/cap_fifo_din_p1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_p1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/cap_fifo_din_p1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[0]~FF  (.D(n1239), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2478)
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp3[0]~FF  (.D(n1240), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp3[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2478)
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp3[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp3[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp3[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp3[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp3[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp3[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp3[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp4[0]~FF  (.D(n1241), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp4[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2478)
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp4[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp4[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp4[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp4[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp4[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp4[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp4[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp5[0]~FF  (.D(n1241), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp5[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2478)
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp5[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp5[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp5[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp5[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp5[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp5[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp5[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp6[0]~FF  (.D(n1240), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp6[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2478)
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp6[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp6[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp6[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp6[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp6[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp6[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp6[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[0]~FF  (.D(n1242), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2478)
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/GEN_PROBE[0].compare_unit_inst/edb_top/la0/tu_data[0]~FF  (.D(n1243), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/tu_data[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2478)
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/edb_top/la0/tu_data[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/edb_top/la0/tu_data[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/edb_top/la0/tu_data[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/edb_top/la0/tu_data[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/edb_top/la0/tu_data[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/edb_top/la0/tu_data[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/edb_top/la0/tu_data[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[1]~FF  (.D(n1244), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2478)
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[2]~FF  (.D(n1245), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2478)
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[3]~FF  (.D(n1246), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2478)
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[4]~FF  (.D(n1247), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2478)
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[5]~FF  (.D(n1248), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2478)
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[6]~FF  (.D(n1249), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2478)
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[7]~FF  (.D(n1250), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2478)
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[1]~FF  (.D(n1251), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2478)
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[2]~FF  (.D(n1252), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2478)
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[3]~FF  (.D(n1253), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2478)
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[4]~FF  (.D(n1254), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2478)
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[5]~FF  (.D(n1255), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2478)
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[6]~FF  (.D(n1256), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2478)
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[7]~FF  (.D(n1257), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2478)
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/trigger_unit_inst/edb_top/la0/tu_trigger~FF  (.D(n1258), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/tu_trigger )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2608)
    defparam \edb_top/la0/trigger_unit_inst/edb_top/la0/tu_trigger~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/trigger_unit_inst/edb_top/la0/tu_trigger~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/trigger_unit_inst/edb_top/la0/tu_trigger~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/trigger_unit_inst/edb_top/la0/tu_trigger~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/trigger_unit_inst/edb_top/la0/tu_trigger~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/trigger_unit_inst/edb_top/la0/tu_trigger~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/trigger_unit_inst/edb_top/la0/tu_trigger~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/cap_fifo_din_cu[1]~FF  (.D(\edb_top/la0/cap_fifo_din_p1[1] ), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/cap_fifo_din_cu[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1649)
    defparam \edb_top/la0/cap_fifo_din_cu[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/cap_fifo_din_cu[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/cap_fifo_din_cu[2]~FF  (.D(\edb_top/la0/cap_fifo_din_p1[2] ), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/cap_fifo_din_cu[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1649)
    defparam \edb_top/la0/cap_fifo_din_cu[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/cap_fifo_din_cu[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/cap_fifo_din_cu[3]~FF  (.D(\edb_top/la0/cap_fifo_din_p1[3] ), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/cap_fifo_din_cu[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1649)
    defparam \edb_top/la0/cap_fifo_din_cu[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/cap_fifo_din_cu[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/cap_fifo_din_cu[4]~FF  (.D(\edb_top/la0/cap_fifo_din_p1[4] ), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/cap_fifo_din_cu[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1649)
    defparam \edb_top/la0/cap_fifo_din_cu[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/cap_fifo_din_cu[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/cap_fifo_din_cu[5]~FF  (.D(\edb_top/la0/cap_fifo_din_p1[5] ), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/cap_fifo_din_cu[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1649)
    defparam \edb_top/la0/cap_fifo_din_cu[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/cap_fifo_din_cu[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/cap_fifo_din_cu[6]~FF  (.D(\edb_top/la0/cap_fifo_din_p1[6] ), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/cap_fifo_din_cu[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1649)
    defparam \edb_top/la0/cap_fifo_din_cu[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/cap_fifo_din_cu[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/cap_fifo_din_cu[7]~FF  (.D(\edb_top/la0/cap_fifo_din_p1[7] ), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/cap_fifo_din_cu[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1649)
    defparam \edb_top/la0/cap_fifo_din_cu[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_cu[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/cap_fifo_din_cu[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/cap_fifo_din_tu[1]~FF  (.D(\edb_top/la0/cap_fifo_din_cu[1] ), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/cap_fifo_din_tu[1]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1661)
    defparam \edb_top/la0/cap_fifo_din_tu[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/cap_fifo_din_tu[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/cap_fifo_din_tu[2]~FF  (.D(\edb_top/la0/cap_fifo_din_cu[2] ), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/cap_fifo_din_tu[2]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1661)
    defparam \edb_top/la0/cap_fifo_din_tu[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/cap_fifo_din_tu[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/cap_fifo_din_tu[3]~FF  (.D(\edb_top/la0/cap_fifo_din_cu[3] ), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/cap_fifo_din_tu[3]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1661)
    defparam \edb_top/la0/cap_fifo_din_tu[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/cap_fifo_din_tu[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/cap_fifo_din_tu[4]~FF  (.D(\edb_top/la0/cap_fifo_din_cu[4] ), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/cap_fifo_din_tu[4]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1661)
    defparam \edb_top/la0/cap_fifo_din_tu[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/cap_fifo_din_tu[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/cap_fifo_din_tu[5]~FF  (.D(\edb_top/la0/cap_fifo_din_cu[5] ), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/cap_fifo_din_tu[5]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1661)
    defparam \edb_top/la0/cap_fifo_din_tu[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/cap_fifo_din_tu[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/cap_fifo_din_tu[6]~FF  (.D(\edb_top/la0/cap_fifo_din_cu[6] ), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/cap_fifo_din_tu[6]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1661)
    defparam \edb_top/la0/cap_fifo_din_tu[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/cap_fifo_din_tu[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/cap_fifo_din_tu[7]~FF  (.D(\edb_top/la0/cap_fifo_din_cu[7] ), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(1'b0), .Q(\edb_top/la0/cap_fifo_din_tu[7]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1661)
    defparam \edb_top/la0/cap_fifo_din_tu[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/cap_fifo_din_tu[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/cap_fifo_din_tu[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/run_trig_p2~FF  (.D(\edb_top/la0/la_biu_inst/run_trig_p1 ), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), .Q(\edb_top/la0/la_biu_inst/run_trig_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1993)
    defparam \edb_top/la0/la_biu_inst/run_trig_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/run_trig_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/run_trig_p2~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/run_trig_p2~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/run_trig_p2~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/run_trig_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/run_trig_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/run_trig_imdt_p1~FF  (.D(\edb_top/la0/la_run_trig_imdt ), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), .Q(\edb_top/la0/la_biu_inst/run_trig_imdt_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1993)
    defparam \edb_top/la0/la_biu_inst/run_trig_imdt_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/run_trig_imdt_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/run_trig_imdt_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/run_trig_imdt_p2~FF  (.D(\edb_top/la0/la_biu_inst/run_trig_imdt_p1 ), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), .Q(\edb_top/la0/la_biu_inst/run_trig_imdt_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1993)
    defparam \edb_top/la0/la_biu_inst/run_trig_imdt_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/run_trig_imdt_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/run_trig_imdt_p2~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/cap_buf_read_done_p1~FF  (.D(n1277), .CE(1'b1), 
           .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), .Q(\edb_top/la0/la_biu_inst/cap_buf_read_done_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1993)
    defparam \edb_top/la0/la_biu_inst/cap_buf_read_done_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/cap_buf_read_done_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/cap_buf_read_done_p1~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/cap_buf_read_done_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/cap_buf_read_done_p1~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/cap_buf_read_done_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/cap_buf_read_done_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/cap_buf_read_done_p2~FF  (.D(\edb_top/la0/la_biu_inst/cap_buf_read_done_p1 ), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), .Q(\edb_top/la0/la_biu_inst/cap_buf_read_done_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1993)
    defparam \edb_top/la0/la_biu_inst/cap_buf_read_done_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/cap_buf_read_done_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/cap_buf_read_done_p2~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/cap_buf_read_done_p2~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/cap_buf_read_done_p2~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/cap_buf_read_done_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/cap_buf_read_done_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/cap_buf_read_done_p3~FF  (.D(\edb_top/la0/la_biu_inst/cap_buf_read_done_p2 ), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), .Q(\edb_top/la0/la_biu_inst/cap_buf_read_done_p3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1993)
    defparam \edb_top/la0/la_biu_inst/cap_buf_read_done_p3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/cap_buf_read_done_p3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/cap_buf_read_done_p3~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/cap_buf_read_done_p3~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/cap_buf_read_done_p3~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/cap_buf_read_done_p3~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/cap_buf_read_done_p3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/pos_counter[12]~FF  (.D(n1282), .CE(n1283), 
           .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), .Q(\edb_top/la0/la_biu_inst/pos_counter[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2014)
    defparam \edb_top/la0/la_biu_inst/pos_counter[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/pos_counter[12]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[12]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/pos_counter[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/edb_top/la0/register_conn[0][0]~FF  (.D(n1284), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), .Q(\edb_top/la0/register_conn[0][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2104)
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/register_conn[0][0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/register_conn[0][0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/register_conn[0][0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/register_conn[0][0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/register_conn[0][0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/register_conn[0][0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/register_conn[0][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/pos_counter[2]~FF  (.D(n1285), .CE(n1283), 
           .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), .Q(\edb_top/la0/la_biu_inst/pos_counter[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2014)
    defparam \edb_top/la0/la_biu_inst/pos_counter[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/pos_counter[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/pos_counter[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/pos_counter[1]~FF  (.D(n1286), .CE(n1283), 
           .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), .Q(\edb_top/la0/la_biu_inst/pos_counter[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2014)
    defparam \edb_top/la0/la_biu_inst/pos_counter[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/pos_counter[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/pos_counter[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/pos_counter[0]~FF  (.D(n1287), .CE(n1283), 
           .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), .Q(\edb_top/la0/la_biu_inst/pos_counter[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2014)
    defparam \edb_top/la0/la_biu_inst/pos_counter[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/pos_counter[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/pos_counter[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/pos_counter[13]~FF  (.D(n1288), .CE(n1283), 
           .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), .Q(\edb_top/la0/la_biu_inst/pos_counter[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2014)
    defparam \edb_top/la0/la_biu_inst/pos_counter[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/pos_counter[13]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[13]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/pos_counter[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/pos_counter[16]~FF  (.D(n1289), .CE(n1283), 
           .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), .Q(\edb_top/la0/la_biu_inst/pos_counter[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2014)
    defparam \edb_top/la0/la_biu_inst/pos_counter[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/pos_counter[16]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[16]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/pos_counter[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/pos_counter[11]~FF  (.D(n1290), .CE(n1283), 
           .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), .Q(\edb_top/la0/la_biu_inst/pos_counter[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2014)
    defparam \edb_top/la0/la_biu_inst/pos_counter[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/pos_counter[11]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[11]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/pos_counter[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/str_sync~FF  (.D(\edb_top/la0/la_biu_inst/str_sync ), 
           .CE(n1292), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_biu_inst/str_sync )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2126)
    defparam \edb_top/la0/la_biu_inst/str_sync~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/str_sync~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/str_sync~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/str_sync~FF .D_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/str_sync~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/str_sync~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/str_sync~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/str_sync_wbff1~FF  (.D(\edb_top/la0/la_biu_inst/str_sync ), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), .Q(\edb_top/la0/la_biu_inst/str_sync_wbff1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2140)
    defparam \edb_top/la0/la_biu_inst/str_sync_wbff1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/str_sync_wbff1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/str_sync_wbff1~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/str_sync_wbff1~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/str_sync_wbff1~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/str_sync_wbff1~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/str_sync_wbff1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/pos_counter[15]~FF  (.D(n1293), .CE(n1283), 
           .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), .Q(\edb_top/la0/la_biu_inst/pos_counter[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2014)
    defparam \edb_top/la0/la_biu_inst/pos_counter[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/pos_counter[15]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[15]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/pos_counter[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/pos_counter[10]~FF  (.D(n1294), .CE(n1283), 
           .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), .Q(\edb_top/la0/la_biu_inst/pos_counter[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2014)
    defparam \edb_top/la0/la_biu_inst/pos_counter[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/pos_counter[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[10]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/pos_counter[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/str_sync_wbff2~FF  (.D(\edb_top/la0/la_biu_inst/str_sync_wbff1 ), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), .Q(\edb_top/la0/la_biu_inst/str_sync_wbff2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2140)
    defparam \edb_top/la0/la_biu_inst/str_sync_wbff2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/str_sync_wbff2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/str_sync_wbff2~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/str_sync_wbff2~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/str_sync_wbff2~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/str_sync_wbff2~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/str_sync_wbff2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/str_sync_wbff2q~FF  (.D(\edb_top/la0/la_biu_inst/str_sync_wbff2 ), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), .Q(\edb_top/la0/la_biu_inst/str_sync_wbff2q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2140)
    defparam \edb_top/la0/la_biu_inst/str_sync_wbff2q~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/str_sync_wbff2q~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/str_sync_wbff2q~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/str_sync_wbff2q~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/str_sync_wbff2q~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/str_sync_wbff2q~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/str_sync_wbff2q~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/rdy_sync~FF  (.D(\edb_top/la0/la_biu_inst/rdy_sync ), 
           .CE(n1298), .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), 
           .Q(\edb_top/la0/la_biu_inst/rdy_sync )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2150)
    defparam \edb_top/la0/la_biu_inst/rdy_sync~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/rdy_sync~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/rdy_sync~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/rdy_sync~FF .D_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/rdy_sync~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/rdy_sync~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/rdy_sync~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/pos_counter[14]~FF  (.D(n1299), .CE(n1283), 
           .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), .Q(\edb_top/la0/la_biu_inst/pos_counter[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2014)
    defparam \edb_top/la0/la_biu_inst/pos_counter[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/pos_counter[14]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[14]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/pos_counter[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/pos_counter[9]~FF  (.D(n1300), .CE(n1283), 
           .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), .Q(\edb_top/la0/la_biu_inst/pos_counter[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2014)
    defparam \edb_top/la0/la_biu_inst/pos_counter[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/pos_counter[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[9]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/pos_counter[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/rdy_sync_tff1~FF  (.D(\edb_top/la0/la_biu_inst/rdy_sync ), 
           .CE(1'b1), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_biu_inst/rdy_sync_tff1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2164)
    defparam \edb_top/la0/la_biu_inst/rdy_sync_tff1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/rdy_sync_tff1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/rdy_sync_tff1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/rdy_sync_tff1~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/rdy_sync_tff1~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/rdy_sync_tff1~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/rdy_sync_tff1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/rdy_sync_tff2~FF  (.D(\edb_top/la0/la_biu_inst/rdy_sync_tff1 ), 
           .CE(1'b1), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_biu_inst/rdy_sync_tff2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2164)
    defparam \edb_top/la0/la_biu_inst/rdy_sync_tff2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/rdy_sync_tff2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/rdy_sync_tff2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/rdy_sync_tff2~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/rdy_sync_tff2~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/rdy_sync_tff2~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/rdy_sync_tff2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/rdy_sync_tff2q~FF  (.D(\edb_top/la0/la_biu_inst/rdy_sync_tff2 ), 
           .CE(1'b1), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_biu_inst/rdy_sync_tff2q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2164)
    defparam \edb_top/la0/la_biu_inst/rdy_sync_tff2q~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/rdy_sync_tff2q~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/rdy_sync_tff2q~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/pos_counter[8]~FF  (.D(n1303), .CE(n1283), 
           .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), .Q(\edb_top/la0/la_biu_inst/pos_counter[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2014)
    defparam \edb_top/la0/la_biu_inst/pos_counter[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/pos_counter[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[8]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/pos_counter[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/pos_counter[7]~FF  (.D(n1304), .CE(n1283), 
           .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), .Q(\edb_top/la0/la_biu_inst/pos_counter[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2014)
    defparam \edb_top/la0/la_biu_inst/pos_counter[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/pos_counter[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[7]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/pos_counter[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/pos_counter[6]~FF  (.D(n1305), .CE(n1283), 
           .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), .Q(\edb_top/la0/la_biu_inst/pos_counter[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2014)
    defparam \edb_top/la0/la_biu_inst/pos_counter[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/pos_counter[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[6]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/pos_counter[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[0]~FF  (.D(\edb_top/la0/la_biu_inst/swapped_data_out[0] ), 
           .CE(n1298), .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), 
           .Q(\edb_top/la0/data_from_biu[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2194)
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/pos_counter[5]~FF  (.D(n1307), .CE(n1283), 
           .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), .Q(\edb_top/la0/la_biu_inst/pos_counter[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2014)
    defparam \edb_top/la0/la_biu_inst/pos_counter[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/pos_counter[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[5]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/pos_counter[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/pos_counter[4]~FF  (.D(n1308), .CE(n1283), 
           .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), .Q(\edb_top/la0/la_biu_inst/pos_counter[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2014)
    defparam \edb_top/la0/la_biu_inst/pos_counter[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/pos_counter[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[4]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/pos_counter[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/axi_fsm_state[0]~FF  (.D(n1309), .CE(n1310), 
           .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), .Q(\edb_top/la0/la_biu_inst/axi_fsm_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2266)
    defparam \edb_top/la0/la_biu_inst/axi_fsm_state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/axi_fsm_state[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/axi_fsm_state[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/pos_counter[3]~FF  (.D(n1311), .CE(n1283), 
           .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), .Q(\edb_top/la0/la_biu_inst/pos_counter[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2014)
    defparam \edb_top/la0/la_biu_inst/pos_counter[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/pos_counter[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[3]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/pos_counter[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/pos_counter[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/run_trig_p1~FF  (.D(\edb_top/la0/la_run_trig ), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), .Q(\edb_top/la0/la_biu_inst/run_trig_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1993)
    defparam \edb_top/la0/la_biu_inst/run_trig_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/run_trig_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/run_trig_p1~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/run_trig_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/run_trig_p1~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/run_trig_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/run_trig_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/edb_top/la0/biu_ready~FF  (.D(n1292), 
           .CE(n1313), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/biu_ready )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2176)
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/biu_ready~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/biu_ready~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/biu_ready~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/biu_ready~FF .D_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/biu_ready~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/biu_ready~FF .SR_VALUE = 1'b1;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/biu_ready~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/edb_top/la0/register_conn[0][1]~FF  (.D(n1314), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), .Q(\edb_top/la0/register_conn[0][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2104)
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/register_conn[0][1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/register_conn[0][1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/register_conn[0][1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/register_conn[0][1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/register_conn[0][1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/register_conn[0][1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/register_conn[0][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/edb_top/la0/register_conn[0][2]~FF  (.D(n1315), 
           .CE(1'b1), .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), .Q(\edb_top/la0/register_conn[0][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2104)
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/register_conn[0][2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/register_conn[0][2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/register_conn[0][2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/register_conn[0][2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/register_conn[0][2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/register_conn[0][2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/register_conn[0][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/row_addr[0]~FF  (.D(\edb_top/la0/address_counter[15] ), 
           .CE(n1292), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_biu_inst/row_addr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2186)
    defparam \edb_top/la0/la_biu_inst/row_addr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/row_addr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/row_addr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/row_addr[1]~FF  (.D(\edb_top/la0/address_counter[16] ), 
           .CE(n1292), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_biu_inst/row_addr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2186)
    defparam \edb_top/la0/la_biu_inst/row_addr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/row_addr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/row_addr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/row_addr[2]~FF  (.D(\edb_top/la0/address_counter[17] ), 
           .CE(n1292), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_biu_inst/row_addr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2186)
    defparam \edb_top/la0/la_biu_inst/row_addr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/row_addr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/row_addr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/row_addr[3]~FF  (.D(\edb_top/la0/address_counter[18] ), 
           .CE(n1292), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_biu_inst/row_addr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2186)
    defparam \edb_top/la0/la_biu_inst/row_addr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/row_addr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/row_addr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/row_addr[4]~FF  (.D(\edb_top/la0/address_counter[19] ), 
           .CE(n1292), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_biu_inst/row_addr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2186)
    defparam \edb_top/la0/la_biu_inst/row_addr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/row_addr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/row_addr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/row_addr[5]~FF  (.D(\edb_top/la0/address_counter[20] ), 
           .CE(n1292), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_biu_inst/row_addr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2186)
    defparam \edb_top/la0/la_biu_inst/row_addr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/row_addr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/row_addr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/row_addr[6]~FF  (.D(\edb_top/la0/address_counter[21] ), 
           .CE(n1292), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_biu_inst/row_addr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2186)
    defparam \edb_top/la0/la_biu_inst/row_addr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/row_addr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/row_addr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/row_addr[7]~FF  (.D(\edb_top/la0/address_counter[22] ), 
           .CE(n1292), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_biu_inst/row_addr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2186)
    defparam \edb_top/la0/la_biu_inst/row_addr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/row_addr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/row_addr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/row_addr[8]~FF  (.D(\edb_top/la0/address_counter[23] ), 
           .CE(n1292), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_biu_inst/row_addr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2186)
    defparam \edb_top/la0/la_biu_inst/row_addr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/row_addr[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/row_addr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/row_addr[9]~FF  (.D(\edb_top/la0/address_counter[24] ), 
           .CE(n1292), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_biu_inst/row_addr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2186)
    defparam \edb_top/la0/la_biu_inst/row_addr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/row_addr[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/row_addr[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/row_addr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[1]~FF  (.D(\edb_top/la0/la_biu_inst/swapped_data_out[1] ), 
           .CE(n1298), .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), 
           .Q(\edb_top/la0/data_from_biu[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2194)
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[2]~FF  (.D(\edb_top/la0/la_biu_inst/swapped_data_out[2] ), 
           .CE(n1298), .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), 
           .Q(\edb_top/la0/data_from_biu[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2194)
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[3]~FF  (.D(\edb_top/la0/la_biu_inst/swapped_data_out[3] ), 
           .CE(n1298), .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), 
           .Q(\edb_top/la0/data_from_biu[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2194)
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[3]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[4]~FF  (.D(\edb_top/la0/la_biu_inst/swapped_data_out[4] ), 
           .CE(n1298), .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), 
           .Q(\edb_top/la0/data_from_biu[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2194)
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[4]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[5]~FF  (.D(\edb_top/la0/la_biu_inst/swapped_data_out[5] ), 
           .CE(n1298), .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), 
           .Q(\edb_top/la0/data_from_biu[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2194)
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[5]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[6]~FF  (.D(\edb_top/la0/la_biu_inst/swapped_data_out[6] ), 
           .CE(n1298), .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), 
           .Q(\edb_top/la0/data_from_biu[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2194)
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[6]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[7]~FF  (.D(\edb_top/la0/la_biu_inst/swapped_data_out[7] ), 
           .CE(n1298), .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), 
           .Q(\edb_top/la0/data_from_biu[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2194)
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[7]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/edb_top/la0/data_from_biu[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/axi_fsm_state[1]~FF  (.D(n1331), .CE(n1310), 
           .CLK(\clk_2~O ), .SR(\edb_top/la0/la_resetn ), .Q(\edb_top/la0/la_biu_inst/axi_fsm_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(2266)
    defparam \edb_top/la0/la_biu_inst/axi_fsm_state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/axi_fsm_state[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/axi_fsm_state[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF  (.D(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0] ), 
           .CE(n1335), .CLK(\clk_2~O ), .SR(n1336), .Q(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1795)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF  (.D(\edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]_2 ), 
           .CE(\edb_top/la0/la_biu_inst/fifo_with_read_inst/we ), .CLK(\clk_2~O ), 
           .SR(n1336), .Q(\edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1786)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF  (.D(n508), 
           .CE(n1335), .CLK(\clk_2~O ), .SR(n1336), .Q(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1795)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF  (.D(n609), 
           .CE(n1335), .CLK(\clk_2~O ), .SR(n1336), .Q(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1795)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF  (.D(n607), 
           .CE(n1335), .CLK(\clk_2~O ), .SR(n1336), .Q(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1795)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF  (.D(n605), 
           .CE(n1335), .CLK(\clk_2~O ), .SR(n1336), .Q(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1795)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF  (.D(n603), 
           .CE(n1335), .CLK(\clk_2~O ), .SR(n1336), .Q(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1795)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF  (.D(n601), 
           .CE(n1335), .CLK(\clk_2~O ), .SR(n1336), .Q(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1795)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF  (.D(n599), 
           .CE(n1335), .CLK(\clk_2~O ), .SR(n1336), .Q(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1795)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF  (.D(n597), 
           .CE(n1335), .CLK(\clk_2~O ), .SR(n1336), .Q(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1795)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF  (.D(n595), 
           .CE(n1335), .CLK(\clk_2~O ), .SR(n1336), .Q(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1795)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF  (.D(n594), 
           .CE(n1335), .CLK(\clk_2~O ), .SR(n1336), .Q(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1795)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF  (.D(n456), 
           .CE(\edb_top/la0/la_biu_inst/fifo_with_read_inst/we ), .CLK(\clk_2~O ), 
           .SR(n1336), .Q(\edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1786)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF  (.D(n626), 
           .CE(\edb_top/la0/la_biu_inst/fifo_with_read_inst/we ), .CLK(\clk_2~O ), 
           .SR(n1336), .Q(\edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1786)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF  (.D(n624), 
           .CE(\edb_top/la0/la_biu_inst/fifo_with_read_inst/we ), .CLK(\clk_2~O ), 
           .SR(n1336), .Q(\edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1786)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF  (.D(n622), 
           .CE(\edb_top/la0/la_biu_inst/fifo_with_read_inst/we ), .CLK(\clk_2~O ), 
           .SR(n1336), .Q(\edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1786)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF  (.D(n620), 
           .CE(\edb_top/la0/la_biu_inst/fifo_with_read_inst/we ), .CLK(\clk_2~O ), 
           .SR(n1336), .Q(\edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1786)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF  (.D(n618), 
           .CE(\edb_top/la0/la_biu_inst/fifo_with_read_inst/we ), .CLK(\clk_2~O ), 
           .SR(n1336), .Q(\edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1786)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF  (.D(n616), 
           .CE(\edb_top/la0/la_biu_inst/fifo_with_read_inst/we ), .CLK(\clk_2~O ), 
           .SR(n1336), .Q(\edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1786)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF  (.D(n614), 
           .CE(\edb_top/la0/la_biu_inst/fifo_with_read_inst/we ), .CLK(\clk_2~O ), 
           .SR(n1336), .Q(\edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1786)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF  (.D(n612), 
           .CE(\edb_top/la0/la_biu_inst/fifo_with_read_inst/we ), .CLK(\clk_2~O ), 
           .SR(n1336), .Q(\edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1786)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF  (.D(n611), 
           .CE(\edb_top/la0/la_biu_inst/fifo_with_read_inst/we ), .CLK(\clk_2~O ), 
           .SR(n1336), .Q(\edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1786)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/internal_register_select[1]~FF  (.D(\edb_top/edb_user_dr[65] ), 
           .CE(n1008), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/internal_register_select[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1036)
    defparam \edb_top/la0/internal_register_select[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/internal_register_select[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/internal_register_select[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/internal_register_select[2]~FF  (.D(\edb_top/edb_user_dr[66] ), 
           .CE(n1008), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/internal_register_select[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1036)
    defparam \edb_top/la0/internal_register_select[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/internal_register_select[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/internal_register_select[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/internal_register_select[3]~FF  (.D(\edb_top/edb_user_dr[67] ), 
           .CE(n1008), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/internal_register_select[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1036)
    defparam \edb_top/la0/internal_register_select[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/internal_register_select[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/internal_register_select[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/internal_register_select[4]~FF  (.D(\edb_top/edb_user_dr[68] ), 
           .CE(n1008), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/internal_register_select[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1036)
    defparam \edb_top/la0/internal_register_select[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/internal_register_select[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/internal_register_select[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/internal_register_select[5]~FF  (.D(\edb_top/edb_user_dr[69] ), 
           .CE(n1008), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/internal_register_select[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1036)
    defparam \edb_top/la0/internal_register_select[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/internal_register_select[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/internal_register_select[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/internal_register_select[6]~FF  (.D(\edb_top/edb_user_dr[70] ), 
           .CE(n1008), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/internal_register_select[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1036)
    defparam \edb_top/la0/internal_register_select[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/internal_register_select[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/internal_register_select[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/internal_register_select[7]~FF  (.D(\edb_top/edb_user_dr[71] ), 
           .CE(n1008), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/internal_register_select[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1036)
    defparam \edb_top/la0/internal_register_select[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/internal_register_select[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/internal_register_select[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/internal_register_select[8]~FF  (.D(\edb_top/edb_user_dr[72] ), 
           .CE(n1008), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/internal_register_select[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1036)
    defparam \edb_top/la0/internal_register_select[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/internal_register_select[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/internal_register_select[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/internal_register_select[9]~FF  (.D(\edb_top/edb_user_dr[73] ), 
           .CE(n1008), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/internal_register_select[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1036)
    defparam \edb_top/la0/internal_register_select[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/internal_register_select[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/internal_register_select[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/internal_register_select[10]~FF  (.D(\edb_top/edb_user_dr[74] ), 
           .CE(n1008), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/internal_register_select[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1036)
    defparam \edb_top/la0/internal_register_select[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/internal_register_select[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/internal_register_select[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/internal_register_select[11]~FF  (.D(\edb_top/edb_user_dr[75] ), 
           .CE(n1008), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/internal_register_select[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1036)
    defparam \edb_top/la0/internal_register_select[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/internal_register_select[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/internal_register_select[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/internal_register_select[12]~FF  (.D(\edb_top/edb_user_dr[76] ), 
           .CE(n1008), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/internal_register_select[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1036)
    defparam \edb_top/la0/internal_register_select[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/internal_register_select[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/internal_register_select[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/internal_register_select[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_pos[1]~FF  (.D(\edb_top/edb_user_dr[46] ), 
           .CE(n978), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_pos[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1073)
    defparam \edb_top/la0/la_trig_pos[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_pos[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_pos[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_pos[2]~FF  (.D(\edb_top/edb_user_dr[47] ), 
           .CE(n978), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_pos[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1073)
    defparam \edb_top/la0/la_trig_pos[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_pos[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_pos[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_pos[3]~FF  (.D(\edb_top/edb_user_dr[48] ), 
           .CE(n978), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_pos[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1073)
    defparam \edb_top/la0/la_trig_pos[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_pos[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_pos[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_pos[4]~FF  (.D(\edb_top/edb_user_dr[49] ), 
           .CE(n978), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_pos[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1073)
    defparam \edb_top/la0/la_trig_pos[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_pos[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_pos[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_pos[5]~FF  (.D(\edb_top/edb_user_dr[50] ), 
           .CE(n978), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_pos[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1073)
    defparam \edb_top/la0/la_trig_pos[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_pos[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_pos[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_pos[6]~FF  (.D(\edb_top/edb_user_dr[51] ), 
           .CE(n978), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_pos[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1073)
    defparam \edb_top/la0/la_trig_pos[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_pos[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_pos[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_pos[7]~FF  (.D(\edb_top/edb_user_dr[52] ), 
           .CE(n978), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_pos[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1073)
    defparam \edb_top/la0/la_trig_pos[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_pos[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_pos[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_pos[8]~FF  (.D(\edb_top/edb_user_dr[53] ), 
           .CE(n978), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_pos[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1073)
    defparam \edb_top/la0/la_trig_pos[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_pos[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_pos[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_pos[9]~FF  (.D(\edb_top/edb_user_dr[54] ), 
           .CE(n978), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_pos[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1073)
    defparam \edb_top/la0/la_trig_pos[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_pos[9]~FF .SR_VALUE = 1'b1;
    defparam \edb_top/la0/la_trig_pos[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_pos[10]~FF  (.D(\edb_top/edb_user_dr[55] ), 
           .CE(n978), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_pos[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1073)
    defparam \edb_top/la0/la_trig_pos[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_pos[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_pos[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_pos[11]~FF  (.D(\edb_top/edb_user_dr[56] ), 
           .CE(n978), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_pos[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1073)
    defparam \edb_top/la0/la_trig_pos[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_pos[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_pos[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_pos[12]~FF  (.D(\edb_top/edb_user_dr[57] ), 
           .CE(n978), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_pos[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1073)
    defparam \edb_top/la0/la_trig_pos[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_pos[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_pos[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_pos[13]~FF  (.D(\edb_top/edb_user_dr[58] ), 
           .CE(n978), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_pos[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1073)
    defparam \edb_top/la0/la_trig_pos[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_pos[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_pos[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_pos[14]~FF  (.D(\edb_top/edb_user_dr[59] ), 
           .CE(n978), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_pos[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1073)
    defparam \edb_top/la0/la_trig_pos[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_pos[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_pos[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_pos[15]~FF  (.D(\edb_top/edb_user_dr[60] ), 
           .CE(n978), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_pos[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1073)
    defparam \edb_top/la0/la_trig_pos[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_pos[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_pos[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/la0/la_trig_pos[16]~FF  (.D(\edb_top/edb_user_dr[61] ), 
           .CE(n978), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/la0/la_trig_pos[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1073)
    defparam \edb_top/la0/la_trig_pos[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/la0/la_trig_pos[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/la0/la_trig_pos[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/la0/la_trig_pos[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/module_id_reg[0]~FF  (.D(\edb_top/edb_user_dr[77] ), 
           .CE(n1514), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/debug_hub_inst/module_id_reg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(307)
    defparam \edb_top/debug_hub_inst/module_id_reg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/module_id_reg[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/module_id_reg[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/module_id_reg[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/module_id_reg[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/module_id_reg[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/module_id_reg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[0]~FF  (.D(\edb_top/edb_user_dr[1] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/module_id_reg[1]~FF  (.D(\edb_top/edb_user_dr[78] ), 
           .CE(n1514), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/debug_hub_inst/module_id_reg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(307)
    defparam \edb_top/debug_hub_inst/module_id_reg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/module_id_reg[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/module_id_reg[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/module_id_reg[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/module_id_reg[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/module_id_reg[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/module_id_reg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/module_id_reg[2]~FF  (.D(\edb_top/edb_user_dr[79] ), 
           .CE(n1514), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/debug_hub_inst/module_id_reg[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(307)
    defparam \edb_top/debug_hub_inst/module_id_reg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/module_id_reg[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/module_id_reg[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/module_id_reg[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/module_id_reg[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/module_id_reg[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/module_id_reg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/module_id_reg[3]~FF  (.D(\edb_top/edb_user_dr[80] ), 
           .CE(n1514), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/debug_hub_inst/module_id_reg[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(307)
    defparam \edb_top/debug_hub_inst/module_id_reg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/module_id_reg[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/module_id_reg[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/module_id_reg[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/module_id_reg[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/module_id_reg[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/module_id_reg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[1]~FF  (.D(\edb_top/edb_user_dr[2] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[2]~FF  (.D(\edb_top/edb_user_dr[3] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[3]~FF  (.D(\edb_top/edb_user_dr[4] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[4]~FF  (.D(\edb_top/edb_user_dr[5] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[5]~FF  (.D(\edb_top/edb_user_dr[6] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[6]~FF  (.D(\edb_top/edb_user_dr[7] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[7]~FF  (.D(\edb_top/edb_user_dr[8] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[8]~FF  (.D(\edb_top/edb_user_dr[9] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[9]~FF  (.D(\edb_top/edb_user_dr[10] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[10]~FF  (.D(\edb_top/edb_user_dr[11] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[11]~FF  (.D(\edb_top/edb_user_dr[12] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[12]~FF  (.D(\edb_top/edb_user_dr[13] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[13]~FF  (.D(\edb_top/edb_user_dr[14] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[14]~FF  (.D(\edb_top/edb_user_dr[15] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[15]~FF  (.D(\edb_top/edb_user_dr[16] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[16]~FF  (.D(\edb_top/edb_user_dr[17] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[17]~FF  (.D(\edb_top/edb_user_dr[18] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[18]~FF  (.D(\edb_top/edb_user_dr[19] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[19]~FF  (.D(\edb_top/edb_user_dr[20] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[20]~FF  (.D(\edb_top/edb_user_dr[21] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[21]~FF  (.D(\edb_top/edb_user_dr[22] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[22]~FF  (.D(\edb_top/edb_user_dr[23] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[23]~FF  (.D(\edb_top/edb_user_dr[24] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[24]~FF  (.D(\edb_top/edb_user_dr[25] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[25]~FF  (.D(\edb_top/edb_user_dr[26] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[26]~FF  (.D(\edb_top/edb_user_dr[27] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[27]~FF  (.D(\edb_top/edb_user_dr[28] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[28]~FF  (.D(\edb_top/edb_user_dr[29] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[29]~FF  (.D(\edb_top/edb_user_dr[30] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[30]~FF  (.D(\edb_top/edb_user_dr[31] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[31]~FF  (.D(\edb_top/edb_user_dr[32] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[32]~FF  (.D(\edb_top/edb_user_dr[33] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[32]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[33]~FF  (.D(\edb_top/edb_user_dr[34] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[33]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[34]~FF  (.D(\edb_top/edb_user_dr[35] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[34]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[35]~FF  (.D(\edb_top/edb_user_dr[36] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[35]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[36]~FF  (.D(\edb_top/edb_user_dr[37] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[36]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[37]~FF  (.D(\edb_top/edb_user_dr[38] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[37]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[38]~FF  (.D(\edb_top/edb_user_dr[39] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[38]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[38]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[39]~FF  (.D(\edb_top/edb_user_dr[40] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[39]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[39]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[40]~FF  (.D(\edb_top/edb_user_dr[41] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[40]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[41]~FF  (.D(\edb_top/edb_user_dr[42] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[41]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[42]~FF  (.D(\edb_top/edb_user_dr[43] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[42]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[43]~FF  (.D(\edb_top/edb_user_dr[44] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[43]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[43]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[44]~FF  (.D(\edb_top/edb_user_dr[45] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[44]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[44]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[45]~FF  (.D(\edb_top/edb_user_dr[46] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[45]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[45]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[46]~FF  (.D(\edb_top/edb_user_dr[47] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[46]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[46]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[47]~FF  (.D(\edb_top/edb_user_dr[48] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[47]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[47]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[48]~FF  (.D(\edb_top/edb_user_dr[49] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[48]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[48]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[49]~FF  (.D(\edb_top/edb_user_dr[50] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[49]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[49]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[50]~FF  (.D(\edb_top/edb_user_dr[51] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[50]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[50]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[51]~FF  (.D(\edb_top/edb_user_dr[52] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[51]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[51]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[52]~FF  (.D(\edb_top/edb_user_dr[53] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[52]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[52]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[53]~FF  (.D(\edb_top/edb_user_dr[54] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[53]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[53]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[54]~FF  (.D(\edb_top/edb_user_dr[55] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[54]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[54]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[55]~FF  (.D(\edb_top/edb_user_dr[56] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[55]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[55]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[56]~FF  (.D(\edb_top/edb_user_dr[57] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[56]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[56]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[57]~FF  (.D(\edb_top/edb_user_dr[58] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[57]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[57]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[58]~FF  (.D(\edb_top/edb_user_dr[59] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[58]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[58]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[59]~FF  (.D(\edb_top/edb_user_dr[60] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[59]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[59]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[60]~FF  (.D(\edb_top/edb_user_dr[61] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[60]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[60]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[61]~FF  (.D(\edb_top/edb_user_dr[62] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[61]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[61]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[62]~FF  (.D(\edb_top/edb_user_dr[63] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[62]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[62]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[63]~FF  (.D(\edb_top/edb_user_dr[64] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[63]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[63]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[64]~FF  (.D(\edb_top/edb_user_dr[65] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[64] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[64]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[64]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[64]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[64]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[64]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[64]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[64]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[65]~FF  (.D(\edb_top/edb_user_dr[66] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[65] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[65]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[65]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[65]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[65]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[65]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[65]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[65]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[66]~FF  (.D(\edb_top/edb_user_dr[67] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[66] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[66]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[66]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[66]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[66]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[66]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[66]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[66]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[67]~FF  (.D(\edb_top/edb_user_dr[68] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[67] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[67]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[67]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[67]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[67]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[67]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[67]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[67]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[68]~FF  (.D(\edb_top/edb_user_dr[69] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[68] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[68]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[68]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[68]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[68]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[68]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[68]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[68]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[69]~FF  (.D(\edb_top/edb_user_dr[70] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[69] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[69]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[69]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[69]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[69]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[69]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[69]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[69]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[70]~FF  (.D(\edb_top/edb_user_dr[71] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[70] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[70]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[70]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[70]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[70]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[70]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[70]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[70]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[71]~FF  (.D(\edb_top/edb_user_dr[72] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[71] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[71]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[71]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[71]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[71]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[71]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[71]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[71]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[72]~FF  (.D(\edb_top/edb_user_dr[73] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[72] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[72]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[72]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[72]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[72]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[72]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[72]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[72]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[73]~FF  (.D(\edb_top/edb_user_dr[74] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[73] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[73]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[73]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[73]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[73]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[73]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[73]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[73]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[74]~FF  (.D(\edb_top/edb_user_dr[75] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[74] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[74]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[74]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[74]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[74]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[74]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[74]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[74]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[75]~FF  (.D(\edb_top/edb_user_dr[76] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[75] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[75]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[75]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[75]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[75]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[75]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[75]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[75]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[76]~FF  (.D(\edb_top/edb_user_dr[77] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[76] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[76]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[76]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[76]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[76]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[76]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[76]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[76]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[77]~FF  (.D(\edb_top/edb_user_dr[78] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[77] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[77]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[77]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[77]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[77]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[77]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[77]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[77]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[78]~FF  (.D(\edb_top/edb_user_dr[79] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[78] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[78]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[78]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[78]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[78]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[78]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[78]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[78]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[79]~FF  (.D(\edb_top/edb_user_dr[80] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[79] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[79]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[79]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[79]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[79]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[79]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[79]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[79]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[80]~FF  (.D(\edb_top/edb_user_dr[81] ), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[80] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[80]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[80]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[80]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[80]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[80]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[80]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[80]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top/debug_hub_inst/edb_top/edb_user_dr[81]~FF  (.D(bscan_TDI), 
           .CE(n1517), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\edb_top/edb_user_dr[81] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(300)
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[81]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[81]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[81]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[81]~FF .D_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[81]~FF .SR_SYNC = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[81]~FF .SR_VALUE = 1'b0;
    defparam \edb_top/debug_hub_inst/edb_top/edb_user_dr[81]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \cnt[1]~FF  (.D(n847), .CE(1'b1), .CLK(\clk_2~O ), .SR(n972), 
           .Q(\cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \cnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \cnt[1]~FF .SR_POLARITY = 1'b1;
    defparam \cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \cnt[1]~FF .SR_SYNC = 1'b1;
    defparam \cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \cnt[2]~FF  (.D(n845), .CE(1'b1), .CLK(\clk_2~O ), .SR(n972), 
           .Q(\cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \cnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \cnt[2]~FF .SR_POLARITY = 1'b1;
    defparam \cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \cnt[2]~FF .SR_SYNC = 1'b1;
    defparam \cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \cnt[3]~FF  (.D(n843), .CE(1'b1), .CLK(\clk_2~O ), .SR(n972), 
           .Q(\cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \cnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \cnt[3]~FF .SR_POLARITY = 1'b1;
    defparam \cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \cnt[3]~FF .SR_SYNC = 1'b1;
    defparam \cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \cnt[4]~FF  (.D(n838), .CE(1'b1), .CLK(\clk_2~O ), .SR(n972), 
           .Q(\cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \cnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \cnt[4]~FF .SR_POLARITY = 1'b1;
    defparam \cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \cnt[4]~FF .SR_SYNC = 1'b1;
    defparam \cnt[4]~FF .SR_VALUE = 1'b0;
    defparam \cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \cnt[5]~FF  (.D(n836), .CE(1'b1), .CLK(\clk_2~O ), .SR(n972), 
           .Q(\cnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \cnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \cnt[5]~FF .SR_POLARITY = 1'b1;
    defparam \cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \cnt[5]~FF .SR_SYNC = 1'b1;
    defparam \cnt[5]~FF .SR_VALUE = 1'b0;
    defparam \cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \cnt[6]~FF  (.D(n834), .CE(1'b1), .CLK(\clk_2~O ), .SR(n972), 
           .Q(\cnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \cnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \cnt[6]~FF .SR_POLARITY = 1'b1;
    defparam \cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \cnt[6]~FF .SR_SYNC = 1'b1;
    defparam \cnt[6]~FF .SR_VALUE = 1'b0;
    defparam \cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \cnt[7]~FF  (.D(n832), .CE(1'b1), .CLK(\clk_2~O ), .SR(n972), 
           .Q(\cnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \cnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \cnt[7]~FF .SR_POLARITY = 1'b1;
    defparam \cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \cnt[7]~FF .SR_SYNC = 1'b1;
    defparam \cnt[7]~FF .SR_VALUE = 1'b0;
    defparam \cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \cnt[8]~FF  (.D(n830), .CE(1'b1), .CLK(\clk_2~O ), .SR(n972), 
           .Q(\cnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \cnt[8]~FF .CE_POLARITY = 1'b1;
    defparam \cnt[8]~FF .SR_POLARITY = 1'b1;
    defparam \cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \cnt[8]~FF .SR_SYNC = 1'b1;
    defparam \cnt[8]~FF .SR_VALUE = 1'b0;
    defparam \cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \cnt[9]~FF  (.D(n828), .CE(1'b1), .CLK(\clk_2~O ), .SR(n972), 
           .Q(\cnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \cnt[9]~FF .CE_POLARITY = 1'b1;
    defparam \cnt[9]~FF .SR_POLARITY = 1'b1;
    defparam \cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \cnt[9]~FF .SR_SYNC = 1'b1;
    defparam \cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \cnt[10]~FF  (.D(n826), .CE(1'b1), .CLK(\clk_2~O ), .SR(n972), 
           .Q(\cnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \cnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \cnt[10]~FF .CE_POLARITY = 1'b1;
    defparam \cnt[10]~FF .SR_POLARITY = 1'b1;
    defparam \cnt[10]~FF .D_POLARITY = 1'b1;
    defparam \cnt[10]~FF .SR_SYNC = 1'b1;
    defparam \cnt[10]~FF .SR_VALUE = 1'b0;
    defparam \cnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \cnt[11]~FF  (.D(n824), .CE(1'b1), .CLK(\clk_2~O ), .SR(n972), 
           .Q(\cnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \cnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \cnt[11]~FF .CE_POLARITY = 1'b1;
    defparam \cnt[11]~FF .SR_POLARITY = 1'b1;
    defparam \cnt[11]~FF .D_POLARITY = 1'b1;
    defparam \cnt[11]~FF .SR_SYNC = 1'b1;
    defparam \cnt[11]~FF .SR_VALUE = 1'b0;
    defparam \cnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \cnt[12]~FF  (.D(n822), .CE(1'b1), .CLK(\clk_2~O ), .SR(n972), 
           .Q(\cnt[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \cnt[12]~FF .CLK_POLARITY = 1'b1;
    defparam \cnt[12]~FF .CE_POLARITY = 1'b1;
    defparam \cnt[12]~FF .SR_POLARITY = 1'b1;
    defparam \cnt[12]~FF .D_POLARITY = 1'b1;
    defparam \cnt[12]~FF .SR_SYNC = 1'b1;
    defparam \cnt[12]~FF .SR_VALUE = 1'b0;
    defparam \cnt[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \cnt[13]~FF  (.D(n820), .CE(1'b1), .CLK(\clk_2~O ), .SR(n972), 
           .Q(\cnt[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \cnt[13]~FF .CLK_POLARITY = 1'b1;
    defparam \cnt[13]~FF .CE_POLARITY = 1'b1;
    defparam \cnt[13]~FF .SR_POLARITY = 1'b1;
    defparam \cnt[13]~FF .D_POLARITY = 1'b1;
    defparam \cnt[13]~FF .SR_SYNC = 1'b1;
    defparam \cnt[13]~FF .SR_VALUE = 1'b0;
    defparam \cnt[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \cnt[14]~FF  (.D(n818), .CE(1'b1), .CLK(\clk_2~O ), .SR(n972), 
           .Q(\cnt[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \cnt[14]~FF .CLK_POLARITY = 1'b1;
    defparam \cnt[14]~FF .CE_POLARITY = 1'b1;
    defparam \cnt[14]~FF .SR_POLARITY = 1'b1;
    defparam \cnt[14]~FF .D_POLARITY = 1'b1;
    defparam \cnt[14]~FF .SR_SYNC = 1'b1;
    defparam \cnt[14]~FF .SR_VALUE = 1'b0;
    defparam \cnt[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \cnt[15]~FF  (.D(n816), .CE(1'b1), .CLK(\clk_2~O ), .SR(n972), 
           .Q(\cnt[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \cnt[15]~FF .CLK_POLARITY = 1'b1;
    defparam \cnt[15]~FF .CE_POLARITY = 1'b1;
    defparam \cnt[15]~FF .SR_POLARITY = 1'b1;
    defparam \cnt[15]~FF .D_POLARITY = 1'b1;
    defparam \cnt[15]~FF .SR_SYNC = 1'b1;
    defparam \cnt[15]~FF .SR_VALUE = 1'b0;
    defparam \cnt[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \cnt[16]~FF  (.D(n814), .CE(1'b1), .CLK(\clk_2~O ), .SR(n972), 
           .Q(\cnt[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \cnt[16]~FF .CLK_POLARITY = 1'b1;
    defparam \cnt[16]~FF .CE_POLARITY = 1'b1;
    defparam \cnt[16]~FF .SR_POLARITY = 1'b1;
    defparam \cnt[16]~FF .D_POLARITY = 1'b1;
    defparam \cnt[16]~FF .SR_SYNC = 1'b1;
    defparam \cnt[16]~FF .SR_VALUE = 1'b0;
    defparam \cnt[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \cnt[17]~FF  (.D(n812), .CE(1'b1), .CLK(\clk_2~O ), .SR(n972), 
           .Q(\cnt[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \cnt[17]~FF .CLK_POLARITY = 1'b1;
    defparam \cnt[17]~FF .CE_POLARITY = 1'b1;
    defparam \cnt[17]~FF .SR_POLARITY = 1'b1;
    defparam \cnt[17]~FF .D_POLARITY = 1'b1;
    defparam \cnt[17]~FF .SR_SYNC = 1'b1;
    defparam \cnt[17]~FF .SR_VALUE = 1'b0;
    defparam \cnt[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \cnt[18]~FF  (.D(n810), .CE(1'b1), .CLK(\clk_2~O ), .SR(n972), 
           .Q(\cnt[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \cnt[18]~FF .CLK_POLARITY = 1'b1;
    defparam \cnt[18]~FF .CE_POLARITY = 1'b1;
    defparam \cnt[18]~FF .SR_POLARITY = 1'b1;
    defparam \cnt[18]~FF .D_POLARITY = 1'b1;
    defparam \cnt[18]~FF .SR_SYNC = 1'b1;
    defparam \cnt[18]~FF .SR_VALUE = 1'b0;
    defparam \cnt[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \cnt[19]~FF  (.D(n808), .CE(1'b1), .CLK(\clk_2~O ), .SR(n972), 
           .Q(\cnt[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \cnt[19]~FF .CLK_POLARITY = 1'b1;
    defparam \cnt[19]~FF .CE_POLARITY = 1'b1;
    defparam \cnt[19]~FF .SR_POLARITY = 1'b1;
    defparam \cnt[19]~FF .D_POLARITY = 1'b1;
    defparam \cnt[19]~FF .SR_SYNC = 1'b1;
    defparam \cnt[19]~FF .SR_VALUE = 1'b0;
    defparam \cnt[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \cnt[20]~FF  (.D(n806), .CE(1'b1), .CLK(\clk_2~O ), .SR(n972), 
           .Q(\cnt[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \cnt[20]~FF .CLK_POLARITY = 1'b1;
    defparam \cnt[20]~FF .CE_POLARITY = 1'b1;
    defparam \cnt[20]~FF .SR_POLARITY = 1'b1;
    defparam \cnt[20]~FF .D_POLARITY = 1'b1;
    defparam \cnt[20]~FF .SR_SYNC = 1'b1;
    defparam \cnt[20]~FF .SR_VALUE = 1'b0;
    defparam \cnt[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \cnt[21]~FF  (.D(n804), .CE(1'b1), .CLK(\clk_2~O ), .SR(n972), 
           .Q(\cnt[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \cnt[21]~FF .CLK_POLARITY = 1'b1;
    defparam \cnt[21]~FF .CE_POLARITY = 1'b1;
    defparam \cnt[21]~FF .SR_POLARITY = 1'b1;
    defparam \cnt[21]~FF .D_POLARITY = 1'b1;
    defparam \cnt[21]~FF .SR_SYNC = 1'b1;
    defparam \cnt[21]~FF .SR_VALUE = 1'b0;
    defparam \cnt[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \cnt[22]~FF  (.D(n802), .CE(1'b1), .CLK(\clk_2~O ), .SR(n972), 
           .Q(\cnt[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \cnt[22]~FF .CLK_POLARITY = 1'b1;
    defparam \cnt[22]~FF .CE_POLARITY = 1'b1;
    defparam \cnt[22]~FF .SR_POLARITY = 1'b1;
    defparam \cnt[22]~FF .D_POLARITY = 1'b1;
    defparam \cnt[22]~FF .SR_SYNC = 1'b1;
    defparam \cnt[22]~FF .SR_VALUE = 1'b0;
    defparam \cnt[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \cnt[23]~FF  (.D(n800), .CE(1'b1), .CLK(\clk_2~O ), .SR(n972), 
           .Q(\cnt[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \cnt[23]~FF .CLK_POLARITY = 1'b1;
    defparam \cnt[23]~FF .CE_POLARITY = 1'b1;
    defparam \cnt[23]~FF .SR_POLARITY = 1'b1;
    defparam \cnt[23]~FF .D_POLARITY = 1'b1;
    defparam \cnt[23]~FF .SR_SYNC = 1'b1;
    defparam \cnt[23]~FF .SR_VALUE = 1'b0;
    defparam \cnt[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \cnt[24]~FF  (.D(n798), .CE(1'b1), .CLK(\clk_2~O ), .SR(n972), 
           .Q(\cnt[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \cnt[24]~FF .CLK_POLARITY = 1'b1;
    defparam \cnt[24]~FF .CE_POLARITY = 1'b1;
    defparam \cnt[24]~FF .SR_POLARITY = 1'b1;
    defparam \cnt[24]~FF .D_POLARITY = 1'b1;
    defparam \cnt[24]~FF .SR_SYNC = 1'b1;
    defparam \cnt[24]~FF .SR_VALUE = 1'b0;
    defparam \cnt[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \cnt[25]~FF  (.D(n796), .CE(1'b1), .CLK(\clk_2~O ), .SR(n972), 
           .Q(\cnt[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \cnt[25]~FF .CLK_POLARITY = 1'b1;
    defparam \cnt[25]~FF .CE_POLARITY = 1'b1;
    defparam \cnt[25]~FF .SR_POLARITY = 1'b1;
    defparam \cnt[25]~FF .D_POLARITY = 1'b1;
    defparam \cnt[25]~FF .SR_SYNC = 1'b1;
    defparam \cnt[25]~FF .SR_VALUE = 1'b0;
    defparam \cnt[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \cnt[26]~FF  (.D(n794), .CE(1'b1), .CLK(\clk_2~O ), .SR(n972), 
           .Q(\cnt[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \cnt[26]~FF .CLK_POLARITY = 1'b1;
    defparam \cnt[26]~FF .CE_POLARITY = 1'b1;
    defparam \cnt[26]~FF .SR_POLARITY = 1'b1;
    defparam \cnt[26]~FF .D_POLARITY = 1'b1;
    defparam \cnt[26]~FF .SR_SYNC = 1'b1;
    defparam \cnt[26]~FF .SR_VALUE = 1'b0;
    defparam \cnt[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \cnt[27]~FF  (.D(n792), .CE(1'b1), .CLK(\clk_2~O ), .SR(n972), 
           .Q(\cnt[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \cnt[27]~FF .CLK_POLARITY = 1'b1;
    defparam \cnt[27]~FF .CE_POLARITY = 1'b1;
    defparam \cnt[27]~FF .SR_POLARITY = 1'b1;
    defparam \cnt[27]~FF .D_POLARITY = 1'b1;
    defparam \cnt[27]~FF .SR_SYNC = 1'b1;
    defparam \cnt[27]~FF .SR_VALUE = 1'b0;
    defparam \cnt[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \cnt[28]~FF  (.D(n790), .CE(1'b1), .CLK(\clk_2~O ), .SR(n972), 
           .Q(\cnt[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \cnt[28]~FF .CLK_POLARITY = 1'b1;
    defparam \cnt[28]~FF .CE_POLARITY = 1'b1;
    defparam \cnt[28]~FF .SR_POLARITY = 1'b1;
    defparam \cnt[28]~FF .D_POLARITY = 1'b1;
    defparam \cnt[28]~FF .SR_SYNC = 1'b1;
    defparam \cnt[28]~FF .SR_VALUE = 1'b0;
    defparam \cnt[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \cnt[29]~FF  (.D(n788), .CE(1'b1), .CLK(\clk_2~O ), .SR(n972), 
           .Q(\cnt[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \cnt[29]~FF .CLK_POLARITY = 1'b1;
    defparam \cnt[29]~FF .CE_POLARITY = 1'b1;
    defparam \cnt[29]~FF .SR_POLARITY = 1'b1;
    defparam \cnt[29]~FF .D_POLARITY = 1'b1;
    defparam \cnt[29]~FF .SR_SYNC = 1'b1;
    defparam \cnt[29]~FF .SR_VALUE = 1'b0;
    defparam \cnt[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \cnt[30]~FF  (.D(n787), .CE(1'b1), .CLK(\clk_2~O ), .SR(n972), 
           .Q(\cnt[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \cnt[30]~FF .CLK_POLARITY = 1'b1;
    defparam \cnt[30]~FF .CE_POLARITY = 1'b1;
    defparam \cnt[30]~FF .SR_POLARITY = 1'b1;
    defparam \cnt[30]~FF .D_POLARITY = 1'b1;
    defparam \cnt[30]~FF .SR_SYNC = 1'b1;
    defparam \cnt[30]~FF .SR_VALUE = 1'b0;
    defparam \cnt[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_ADD \edb_top/la0/add_45/i2  (.I0(\edb_top/la0/address_counter[16] ), 
            .I1(\edb_top/la0/address_counter[15] ), .CI(1'b0), .O(n24), 
            .CO(n25)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1092)
    defparam \edb_top/la0/add_45/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_45/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_46/i1  (.I0(\edb_top/la0/address_counter[0] ), 
            .I1(n986), .CI(1'b0), .O(n34), .CO(n35)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1093)
    defparam \edb_top/la0/add_46/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_46/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_52/i2  (.I0(\edb_top/la0/bit_count[1] ), .I1(\edb_top/la0/bit_count[0] ), 
            .CI(1'b0), .O(n36), .CO(n37)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1120)
    defparam \edb_top/la0/add_52/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_52/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/sub_59/add_2/i1  (.I0(\edb_top/la0/word_count[0] ), 
            .I1(1'b0), .CI(n2038), .O(n40), .CO(n41)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1130)
    defparam \edb_top/la0/sub_59/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/sub_59/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_13/i2  (.I0(\edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]_2 ), 
            .I1(\edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]_2 ), 
            .CI(1'b0), .O(n456), .CO(n457)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1784)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_13/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_13/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_18/i2  (.I0(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1] ), 
            .I1(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0] ), 
            .CI(1'b0), .O(n508), .CO(n509)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1793)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_18/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_18/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_22/i1  (.I0(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0] ), 
            .I1(\edb_top/la0/la_biu_inst/row_addr[0] ), .CI(1'b0), .O(n511), 
            .CO(n512)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1797)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_22/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_22/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/debug_hub_inst/sub_28/add_2/i1  (.I0(\edb_top/debug_hub_inst/module_id_reg[0] ), 
            .I1(1'b0), .CI(n2039), .O(n532), .CO(n533)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(324)
    defparam \edb_top/debug_hub_inst/sub_28/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/sub_28/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/debug_hub_inst/sub_28/add_2/i2  (.I0(\edb_top/debug_hub_inst/module_id_reg[1] ), 
            .I1(1'b1), .CI(n533), .O(n534), .CO(n535)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(324)
    defparam \edb_top/debug_hub_inst/sub_28/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/sub_28/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/debug_hub_inst/sub_28/add_2/i4  (.I0(\edb_top/debug_hub_inst/module_id_reg[3] ), 
            .I1(1'b1), .CI(n576), .O(n574)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(324)
    defparam \edb_top/debug_hub_inst/sub_28/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/sub_28/add_2/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/debug_hub_inst/sub_28/add_2/i3  (.I0(\edb_top/debug_hub_inst/module_id_reg[2] ), 
            .I1(1'b1), .CI(n535), .O(n575), .CO(n576)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(324)
    defparam \edb_top/debug_hub_inst/sub_28/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top/debug_hub_inst/sub_28/add_2/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_22/i10  (.I0(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9] ), 
            .I1(\edb_top/la0/la_biu_inst/row_addr[9] ), .CI(n579), .O(n577)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1797)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_22/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_22/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_22/i9  (.I0(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8] ), 
            .I1(\edb_top/la0/la_biu_inst/row_addr[8] ), .CI(n581), .O(n578), 
            .CO(n579)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1797)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_22/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_22/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_22/i8  (.I0(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7] ), 
            .I1(\edb_top/la0/la_biu_inst/row_addr[7] ), .CI(n583), .O(n580), 
            .CO(n581)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1797)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_22/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_22/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_22/i7  (.I0(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6] ), 
            .I1(\edb_top/la0/la_biu_inst/row_addr[6] ), .CI(n585), .O(n582), 
            .CO(n583)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1797)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_22/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_22/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_22/i6  (.I0(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5] ), 
            .I1(\edb_top/la0/la_biu_inst/row_addr[5] ), .CI(n587), .O(n584), 
            .CO(n585)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1797)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_22/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_22/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_22/i5  (.I0(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4] ), 
            .I1(\edb_top/la0/la_biu_inst/row_addr[4] ), .CI(n589), .O(n586), 
            .CO(n587)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1797)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_22/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_22/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_22/i4  (.I0(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3] ), 
            .I1(\edb_top/la0/la_biu_inst/row_addr[3] ), .CI(n591), .O(n588), 
            .CO(n589)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1797)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_22/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_22/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_22/i3  (.I0(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2] ), 
            .I1(\edb_top/la0/la_biu_inst/row_addr[2] ), .CI(n593), .O(n590), 
            .CO(n591)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1797)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_22/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_22/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_22/i2  (.I0(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1] ), 
            .I1(\edb_top/la0/la_biu_inst/row_addr[1] ), .CI(n512), .O(n592), 
            .CO(n593)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1797)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_22/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_22/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_18/i11  (.I0(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10] ), 
            .I1(1'b0), .CI(n596), .O(n594)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1793)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_18/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_18/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_18/i10  (.I0(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9] ), 
            .I1(1'b0), .CI(n598), .O(n595), .CO(n596)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1793)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_18/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_18/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_18/i9  (.I0(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8] ), 
            .I1(1'b0), .CI(n600), .O(n597), .CO(n598)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1793)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_18/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_18/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_18/i8  (.I0(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7] ), 
            .I1(1'b0), .CI(n602), .O(n599), .CO(n600)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1793)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_18/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_18/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_18/i7  (.I0(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6] ), 
            .I1(1'b0), .CI(n604), .O(n601), .CO(n602)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1793)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_18/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_18/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_18/i6  (.I0(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5] ), 
            .I1(1'b0), .CI(n606), .O(n603), .CO(n604)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1793)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_18/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_18/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_18/i5  (.I0(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4] ), 
            .I1(1'b0), .CI(n608), .O(n605), .CO(n606)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1793)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_18/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_18/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_18/i4  (.I0(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3] ), 
            .I1(1'b0), .CI(n610), .O(n607), .CO(n608)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1793)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_18/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_18/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_18/i3  (.I0(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2] ), 
            .I1(1'b0), .CI(n509), .O(n609), .CO(n610)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1793)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_18/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_18/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_13/i11  (.I0(\edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] ), 
            .I1(1'b0), .CI(n613), .O(n611)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1784)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_13/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_13/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_13/i10  (.I0(\edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]_2 ), 
            .I1(1'b0), .CI(n615), .O(n612), .CO(n613)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1784)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_13/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_13/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_13/i9  (.I0(\edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]_2 ), 
            .I1(1'b0), .CI(n617), .O(n614), .CO(n615)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1784)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_13/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_13/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_13/i8  (.I0(\edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]_2 ), 
            .I1(1'b0), .CI(n619), .O(n616), .CO(n617)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1784)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_13/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_13/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_13/i7  (.I0(\edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]_2 ), 
            .I1(1'b0), .CI(n621), .O(n618), .CO(n619)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1784)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_13/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_13/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_13/i6  (.I0(\edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]_2 ), 
            .I1(1'b0), .CI(n623), .O(n620), .CO(n621)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1784)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_13/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_13/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_13/i5  (.I0(\edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]_2 ), 
            .I1(1'b0), .CI(n625), .O(n622), .CO(n623)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1784)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_13/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_13/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_13/i4  (.I0(\edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]_2 ), 
            .I1(1'b0), .CI(n627), .O(n624), .CO(n625)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1784)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_13/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_13/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_13/i3  (.I0(\edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]_2 ), 
            .I1(1'b0), .CI(n457), .O(n626), .CO(n627)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1784)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_13/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/add_13/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/add_12/i17  (.I0(\edb_top/la0/la_biu_inst/pos_counter[16] ), 
            .I1(1'b0), .CI(n630), .O(n628)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1996)
    defparam \edb_top/la0/la_biu_inst/add_12/i17 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/add_12/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/add_12/i16  (.I0(\edb_top/la0/la_biu_inst/pos_counter[15] ), 
            .I1(1'b0), .CI(n632), .O(n629), .CO(n630)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1996)
    defparam \edb_top/la0/la_biu_inst/add_12/i16 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/add_12/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/add_12/i15  (.I0(\edb_top/la0/la_biu_inst/pos_counter[14] ), 
            .I1(1'b0), .CI(n634), .O(n631), .CO(n632)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1996)
    defparam \edb_top/la0/la_biu_inst/add_12/i15 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/add_12/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/add_12/i14  (.I0(\edb_top/la0/la_biu_inst/pos_counter[13] ), 
            .I1(1'b0), .CI(n636), .O(n633), .CO(n634)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1996)
    defparam \edb_top/la0/la_biu_inst/add_12/i14 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/add_12/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/add_12/i13  (.I0(\edb_top/la0/la_biu_inst/pos_counter[12] ), 
            .I1(1'b0), .CI(n638), .O(n635), .CO(n636)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1996)
    defparam \edb_top/la0/la_biu_inst/add_12/i13 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/add_12/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/add_12/i12  (.I0(\edb_top/la0/la_biu_inst/pos_counter[11] ), 
            .I1(1'b0), .CI(n640), .O(n637), .CO(n638)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1996)
    defparam \edb_top/la0/la_biu_inst/add_12/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/add_12/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/add_12/i11  (.I0(\edb_top/la0/la_biu_inst/pos_counter[10] ), 
            .I1(1'b0), .CI(n642), .O(n639), .CO(n640)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1996)
    defparam \edb_top/la0/la_biu_inst/add_12/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/add_12/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/add_12/i10  (.I0(\edb_top/la0/la_biu_inst/pos_counter[9] ), 
            .I1(1'b0), .CI(n644), .O(n641), .CO(n642)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1996)
    defparam \edb_top/la0/la_biu_inst/add_12/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/add_12/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/add_12/i9  (.I0(\edb_top/la0/la_biu_inst/pos_counter[8] ), 
            .I1(1'b0), .CI(n646), .O(n643), .CO(n644)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1996)
    defparam \edb_top/la0/la_biu_inst/add_12/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/add_12/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/add_12/i8  (.I0(\edb_top/la0/la_biu_inst/pos_counter[7] ), 
            .I1(1'b0), .CI(n648), .O(n645), .CO(n646)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1996)
    defparam \edb_top/la0/la_biu_inst/add_12/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/add_12/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/add_12/i7  (.I0(\edb_top/la0/la_biu_inst/pos_counter[6] ), 
            .I1(1'b0), .CI(n650), .O(n647), .CO(n648)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1996)
    defparam \edb_top/la0/la_biu_inst/add_12/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/add_12/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/add_12/i6  (.I0(\edb_top/la0/la_biu_inst/pos_counter[5] ), 
            .I1(1'b0), .CI(n652), .O(n649), .CO(n650)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1996)
    defparam \edb_top/la0/la_biu_inst/add_12/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/add_12/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/add_12/i5  (.I0(\edb_top/la0/la_biu_inst/pos_counter[4] ), 
            .I1(1'b0), .CI(n654), .O(n651), .CO(n652)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1996)
    defparam \edb_top/la0/la_biu_inst/add_12/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/add_12/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/add_12/i4  (.I0(\edb_top/la0/la_biu_inst/pos_counter[3] ), 
            .I1(1'b0), .CI(n656), .O(n653), .CO(n654)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1996)
    defparam \edb_top/la0/la_biu_inst/add_12/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/add_12/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/add_12/i3  (.I0(\edb_top/la0/la_biu_inst/pos_counter[2] ), 
            .I1(1'b0), .CI(n658), .O(n655), .CO(n656)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1996)
    defparam \edb_top/la0/la_biu_inst/add_12/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/add_12/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/la_biu_inst/add_12/i2  (.I0(\edb_top/la0/la_biu_inst/pos_counter[1] ), 
            .I1(\edb_top/la0/la_biu_inst/pos_counter[0] ), .CI(1'b0), .O(n657), 
            .CO(n658)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1996)
    defparam \edb_top/la0/la_biu_inst/add_12/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/add_12/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/sub_59/add_2/i16  (.I0(\edb_top/la0/word_count[15] ), 
            .I1(1'b1), .CI(n661), .O(n659)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1130)
    defparam \edb_top/la0/sub_59/add_2/i16 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/sub_59/add_2/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/sub_59/add_2/i15  (.I0(\edb_top/la0/word_count[14] ), 
            .I1(1'b1), .CI(n663), .O(n660), .CO(n661)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1130)
    defparam \edb_top/la0/sub_59/add_2/i15 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/sub_59/add_2/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/sub_59/add_2/i14  (.I0(\edb_top/la0/word_count[13] ), 
            .I1(1'b1), .CI(n665), .O(n662), .CO(n663)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1130)
    defparam \edb_top/la0/sub_59/add_2/i14 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/sub_59/add_2/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/sub_59/add_2/i13  (.I0(\edb_top/la0/word_count[12] ), 
            .I1(1'b1), .CI(n667), .O(n664), .CO(n665)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1130)
    defparam \edb_top/la0/sub_59/add_2/i13 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/sub_59/add_2/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/sub_59/add_2/i12  (.I0(\edb_top/la0/word_count[11] ), 
            .I1(1'b1), .CI(n669), .O(n666), .CO(n667)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1130)
    defparam \edb_top/la0/sub_59/add_2/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/sub_59/add_2/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/sub_59/add_2/i11  (.I0(\edb_top/la0/word_count[10] ), 
            .I1(1'b1), .CI(n671), .O(n668), .CO(n669)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1130)
    defparam \edb_top/la0/sub_59/add_2/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/sub_59/add_2/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/sub_59/add_2/i10  (.I0(\edb_top/la0/word_count[9] ), 
            .I1(1'b1), .CI(n673), .O(n670), .CO(n671)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1130)
    defparam \edb_top/la0/sub_59/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/sub_59/add_2/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/sub_59/add_2/i9  (.I0(\edb_top/la0/word_count[8] ), 
            .I1(1'b1), .CI(n675), .O(n672), .CO(n673)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1130)
    defparam \edb_top/la0/sub_59/add_2/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/sub_59/add_2/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/sub_59/add_2/i8  (.I0(\edb_top/la0/word_count[7] ), 
            .I1(1'b1), .CI(n677), .O(n674), .CO(n675)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1130)
    defparam \edb_top/la0/sub_59/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/sub_59/add_2/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/sub_59/add_2/i7  (.I0(\edb_top/la0/word_count[6] ), 
            .I1(1'b1), .CI(n679), .O(n676), .CO(n677)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1130)
    defparam \edb_top/la0/sub_59/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/sub_59/add_2/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/sub_59/add_2/i6  (.I0(\edb_top/la0/word_count[5] ), 
            .I1(1'b1), .CI(n681), .O(n678), .CO(n679)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1130)
    defparam \edb_top/la0/sub_59/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/sub_59/add_2/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/sub_59/add_2/i5  (.I0(\edb_top/la0/word_count[4] ), 
            .I1(1'b1), .CI(n683), .O(n680), .CO(n681)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1130)
    defparam \edb_top/la0/sub_59/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/sub_59/add_2/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/sub_59/add_2/i4  (.I0(\edb_top/la0/word_count[3] ), 
            .I1(1'b1), .CI(n685), .O(n682), .CO(n683)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1130)
    defparam \edb_top/la0/sub_59/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/sub_59/add_2/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/sub_59/add_2/i3  (.I0(\edb_top/la0/word_count[2] ), 
            .I1(1'b1), .CI(n687), .O(n684), .CO(n685)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1130)
    defparam \edb_top/la0/sub_59/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/sub_59/add_2/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/sub_59/add_2/i2  (.I0(\edb_top/la0/word_count[1] ), 
            .I1(1'b1), .CI(n41), .O(n686), .CO(n687)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1130)
    defparam \edb_top/la0/sub_59/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/sub_59/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_52/i6  (.I0(\edb_top/la0/bit_count[5] ), .I1(1'b0), 
            .CI(n692), .O(n689)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1120)
    defparam \edb_top/la0/add_52/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_52/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_52/i5  (.I0(\edb_top/la0/bit_count[4] ), .I1(1'b0), 
            .CI(n694), .O(n691), .CO(n692)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1120)
    defparam \edb_top/la0/add_52/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_52/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_52/i4  (.I0(\edb_top/la0/bit_count[3] ), .I1(1'b0), 
            .CI(n696), .O(n693), .CO(n694)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1120)
    defparam \edb_top/la0/add_52/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_52/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_52/i3  (.I0(\edb_top/la0/bit_count[2] ), .I1(1'b0), 
            .CI(n37), .O(n695), .CO(n696)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1120)
    defparam \edb_top/la0/add_52/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_52/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_46/i25  (.I0(\edb_top/la0/address_counter[24] ), 
            .I1(1'b0), .CI(n713), .O(n710)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1093)
    defparam \edb_top/la0/add_46/i25 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_46/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_46/i24  (.I0(\edb_top/la0/address_counter[23] ), 
            .I1(1'b0), .CI(n715), .O(n712), .CO(n713)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1093)
    defparam \edb_top/la0/add_46/i24 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_46/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_46/i23  (.I0(\edb_top/la0/address_counter[22] ), 
            .I1(1'b0), .CI(n717), .O(n714), .CO(n715)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1093)
    defparam \edb_top/la0/add_46/i23 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_46/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_46/i22  (.I0(\edb_top/la0/address_counter[21] ), 
            .I1(1'b0), .CI(n719), .O(n716), .CO(n717)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1093)
    defparam \edb_top/la0/add_46/i22 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_46/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_46/i21  (.I0(\edb_top/la0/address_counter[20] ), 
            .I1(1'b0), .CI(n721), .O(n718), .CO(n719)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1093)
    defparam \edb_top/la0/add_46/i21 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_46/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_46/i20  (.I0(\edb_top/la0/address_counter[19] ), 
            .I1(1'b0), .CI(n723), .O(n720), .CO(n721)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1093)
    defparam \edb_top/la0/add_46/i20 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_46/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_46/i19  (.I0(\edb_top/la0/address_counter[18] ), 
            .I1(1'b0), .CI(n725), .O(n722), .CO(n723)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1093)
    defparam \edb_top/la0/add_46/i19 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_46/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_46/i18  (.I0(\edb_top/la0/address_counter[17] ), 
            .I1(1'b0), .CI(n727), .O(n724), .CO(n725)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1093)
    defparam \edb_top/la0/add_46/i18 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_46/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_46/i17  (.I0(\edb_top/la0/address_counter[16] ), 
            .I1(1'b0), .CI(n729), .O(n726), .CO(n727)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1093)
    defparam \edb_top/la0/add_46/i17 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_46/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_46/i16  (.I0(\edb_top/la0/address_counter[15] ), 
            .I1(1'b0), .CI(n731), .O(n728), .CO(n729)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1093)
    defparam \edb_top/la0/add_46/i16 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_46/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_46/i15  (.I0(\edb_top/la0/address_counter[14] ), 
            .I1(1'b0), .CI(n733), .O(n730), .CO(n731)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1093)
    defparam \edb_top/la0/add_46/i15 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_46/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_46/i14  (.I0(\edb_top/la0/address_counter[13] ), 
            .I1(1'b0), .CI(n735), .O(n732), .CO(n733)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1093)
    defparam \edb_top/la0/add_46/i14 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_46/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_46/i13  (.I0(\edb_top/la0/address_counter[12] ), 
            .I1(1'b0), .CI(n737), .O(n734), .CO(n735)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1093)
    defparam \edb_top/la0/add_46/i13 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_46/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_46/i12  (.I0(\edb_top/la0/address_counter[11] ), 
            .I1(1'b0), .CI(n739), .O(n736), .CO(n737)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1093)
    defparam \edb_top/la0/add_46/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_46/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_46/i11  (.I0(\edb_top/la0/address_counter[10] ), 
            .I1(1'b0), .CI(n741), .O(n738), .CO(n739)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1093)
    defparam \edb_top/la0/add_46/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_46/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_46/i10  (.I0(\edb_top/la0/address_counter[9] ), 
            .I1(1'b0), .CI(n743), .O(n740), .CO(n741)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1093)
    defparam \edb_top/la0/add_46/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_46/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_46/i9  (.I0(\edb_top/la0/address_counter[8] ), 
            .I1(1'b0), .CI(n745), .O(n742), .CO(n743)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1093)
    defparam \edb_top/la0/add_46/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_46/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_46/i8  (.I0(\edb_top/la0/address_counter[7] ), 
            .I1(1'b0), .CI(n747), .O(n744), .CO(n745)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1093)
    defparam \edb_top/la0/add_46/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_46/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_46/i7  (.I0(\edb_top/la0/address_counter[6] ), 
            .I1(1'b0), .CI(n749), .O(n746), .CO(n747)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1093)
    defparam \edb_top/la0/add_46/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_46/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_46/i6  (.I0(\edb_top/la0/address_counter[5] ), 
            .I1(1'b0), .CI(n751), .O(n748), .CO(n749)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1093)
    defparam \edb_top/la0/add_46/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_46/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_46/i5  (.I0(\edb_top/la0/address_counter[4] ), 
            .I1(1'b0), .CI(n753), .O(n750), .CO(n751)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1093)
    defparam \edb_top/la0/add_46/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_46/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_46/i4  (.I0(\edb_top/la0/address_counter[3] ), 
            .I1(1'b0), .CI(n755), .O(n752), .CO(n753)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1093)
    defparam \edb_top/la0/add_46/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_46/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_46/i3  (.I0(\edb_top/la0/address_counter[2] ), 
            .I1(1'b0), .CI(n757), .O(n754), .CO(n755)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1093)
    defparam \edb_top/la0/add_46/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_46/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_46/i2  (.I0(\edb_top/la0/address_counter[1] ), 
            .I1(1'b0), .CI(n35), .O(n756), .CO(n757)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1093)
    defparam \edb_top/la0/add_46/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_46/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_45/i10  (.I0(\edb_top/la0/address_counter[24] ), 
            .I1(1'b0), .CI(n774), .O(n771)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1092)
    defparam \edb_top/la0/add_45/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_45/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_45/i9  (.I0(\edb_top/la0/address_counter[23] ), 
            .I1(1'b0), .CI(n776), .O(n773), .CO(n774)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1092)
    defparam \edb_top/la0/add_45/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_45/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_45/i8  (.I0(\edb_top/la0/address_counter[22] ), 
            .I1(1'b0), .CI(n778), .O(n775), .CO(n776)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1092)
    defparam \edb_top/la0/add_45/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_45/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_45/i7  (.I0(\edb_top/la0/address_counter[21] ), 
            .I1(1'b0), .CI(n780), .O(n777), .CO(n778)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1092)
    defparam \edb_top/la0/add_45/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_45/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_45/i6  (.I0(\edb_top/la0/address_counter[20] ), 
            .I1(1'b0), .CI(n782), .O(n779), .CO(n780)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1092)
    defparam \edb_top/la0/add_45/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_45/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_45/i5  (.I0(\edb_top/la0/address_counter[19] ), 
            .I1(1'b0), .CI(n784), .O(n781), .CO(n782)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1092)
    defparam \edb_top/la0/add_45/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_45/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_45/i4  (.I0(\edb_top/la0/address_counter[18] ), 
            .I1(1'b0), .CI(n786), .O(n783), .CO(n784)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1092)
    defparam \edb_top/la0/add_45/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_45/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top/la0/add_45/i3  (.I0(\edb_top/la0/address_counter[17] ), 
            .I1(1'b0), .CI(n25), .O(n785), .CO(n786)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(1092)
    defparam \edb_top/la0/add_45/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top/la0/add_45/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \add_6/i31  (.I0(\cnt[30] ), .I1(1'b0), .CI(n789), .O(n787)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \add_6/i31 .I0_POLARITY = 1'b1;
    defparam \add_6/i31 .I1_POLARITY = 1'b1;
    EFX_ADD \add_6/i30  (.I0(\cnt[29] ), .I1(1'b0), .CI(n791), .O(n788), 
            .CO(n789)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \add_6/i30 .I0_POLARITY = 1'b1;
    defparam \add_6/i30 .I1_POLARITY = 1'b1;
    EFX_ADD \add_6/i29  (.I0(\cnt[28] ), .I1(1'b0), .CI(n793), .O(n790), 
            .CO(n791)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \add_6/i29 .I0_POLARITY = 1'b1;
    defparam \add_6/i29 .I1_POLARITY = 1'b1;
    EFX_ADD \add_6/i28  (.I0(\cnt[27] ), .I1(1'b0), .CI(n795), .O(n792), 
            .CO(n793)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \add_6/i28 .I0_POLARITY = 1'b1;
    defparam \add_6/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \add_6/i27  (.I0(\cnt[26] ), .I1(1'b0), .CI(n797), .O(n794), 
            .CO(n795)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \add_6/i27 .I0_POLARITY = 1'b1;
    defparam \add_6/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \add_6/i26  (.I0(\cnt[25] ), .I1(1'b0), .CI(n799), .O(n796), 
            .CO(n797)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \add_6/i26 .I0_POLARITY = 1'b1;
    defparam \add_6/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \add_6/i25  (.I0(\cnt[24] ), .I1(1'b0), .CI(n801), .O(n798), 
            .CO(n799)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \add_6/i25 .I0_POLARITY = 1'b1;
    defparam \add_6/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \add_6/i24  (.I0(\cnt[23] ), .I1(1'b0), .CI(n803), .O(n800), 
            .CO(n801)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \add_6/i24 .I0_POLARITY = 1'b1;
    defparam \add_6/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \add_6/i23  (.I0(\cnt[22] ), .I1(1'b0), .CI(n805), .O(n802), 
            .CO(n803)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \add_6/i23 .I0_POLARITY = 1'b1;
    defparam \add_6/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \add_6/i22  (.I0(\cnt[21] ), .I1(1'b0), .CI(n807), .O(n804), 
            .CO(n805)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \add_6/i22 .I0_POLARITY = 1'b1;
    defparam \add_6/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \add_6/i21  (.I0(\cnt[20] ), .I1(1'b0), .CI(n809), .O(n806), 
            .CO(n807)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \add_6/i21 .I0_POLARITY = 1'b1;
    defparam \add_6/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \add_6/i20  (.I0(\cnt[19] ), .I1(1'b0), .CI(n811), .O(n808), 
            .CO(n809)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \add_6/i20 .I0_POLARITY = 1'b1;
    defparam \add_6/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \add_6/i19  (.I0(\cnt[18] ), .I1(1'b0), .CI(n813), .O(n810), 
            .CO(n811)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \add_6/i19 .I0_POLARITY = 1'b1;
    defparam \add_6/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \add_6/i18  (.I0(\cnt[17] ), .I1(1'b0), .CI(n815), .O(n812), 
            .CO(n813)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \add_6/i18 .I0_POLARITY = 1'b1;
    defparam \add_6/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \add_6/i17  (.I0(\cnt[16] ), .I1(1'b0), .CI(n817), .O(n814), 
            .CO(n815)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \add_6/i17 .I0_POLARITY = 1'b1;
    defparam \add_6/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \add_6/i16  (.I0(\cnt[15] ), .I1(1'b0), .CI(n819), .O(n816), 
            .CO(n817)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \add_6/i16 .I0_POLARITY = 1'b1;
    defparam \add_6/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \add_6/i15  (.I0(\cnt[14] ), .I1(1'b0), .CI(n821), .O(n818), 
            .CO(n819)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \add_6/i15 .I0_POLARITY = 1'b1;
    defparam \add_6/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \add_6/i14  (.I0(\cnt[13] ), .I1(1'b0), .CI(n823), .O(n820), 
            .CO(n821)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \add_6/i14 .I0_POLARITY = 1'b1;
    defparam \add_6/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \add_6/i13  (.I0(\cnt[12] ), .I1(1'b0), .CI(n825), .O(n822), 
            .CO(n823)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \add_6/i13 .I0_POLARITY = 1'b1;
    defparam \add_6/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \add_6/i12  (.I0(\cnt[11] ), .I1(1'b0), .CI(n827), .O(n824), 
            .CO(n825)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \add_6/i12 .I0_POLARITY = 1'b1;
    defparam \add_6/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \add_6/i11  (.I0(\cnt[10] ), .I1(1'b0), .CI(n829), .O(n826), 
            .CO(n827)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \add_6/i11 .I0_POLARITY = 1'b1;
    defparam \add_6/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \add_6/i10  (.I0(\cnt[9] ), .I1(1'b0), .CI(n831), .O(n828), 
            .CO(n829)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \add_6/i10 .I0_POLARITY = 1'b1;
    defparam \add_6/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \add_6/i9  (.I0(\cnt[8] ), .I1(1'b0), .CI(n833), .O(n830), 
            .CO(n831)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \add_6/i9 .I0_POLARITY = 1'b1;
    defparam \add_6/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \add_6/i8  (.I0(\cnt[7] ), .I1(1'b0), .CI(n835), .O(n832), 
            .CO(n833)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \add_6/i8 .I0_POLARITY = 1'b1;
    defparam \add_6/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \add_6/i7  (.I0(\cnt[6] ), .I1(1'b0), .CI(n837), .O(n834), 
            .CO(n835)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \add_6/i7 .I0_POLARITY = 1'b1;
    defparam \add_6/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \add_6/i6  (.I0(\cnt[5] ), .I1(1'b0), .CI(n839), .O(n836), 
            .CO(n837)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \add_6/i6 .I0_POLARITY = 1'b1;
    defparam \add_6/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \add_6/i5  (.I0(\cnt[4] ), .I1(1'b0), .CI(n844), .O(n838), 
            .CO(n839)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \add_6/i5 .I0_POLARITY = 1'b1;
    defparam \add_6/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \add_6/i4  (.I0(\cnt[3] ), .I1(1'b0), .CI(n846), .O(n843), 
            .CO(n844)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \add_6/i4 .I0_POLARITY = 1'b1;
    defparam \add_6/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \add_6/i3  (.I0(\cnt[2] ), .I1(1'b0), .CI(n848), .O(n845), 
            .CO(n846)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \add_6/i3 .I0_POLARITY = 1'b1;
    defparam \add_6/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \add_6/i2  (.I0(\cnt[1] ), .I1(\cnt[0] ), .CI(1'b0), .O(n847), 
            .CO(n848)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/top.v(57)
    defparam \add_6/i2 .I0_POLARITY = 1'b1;
    defparam \add_6/i2 .I1_POLARITY = 1'b1;
    EFX_RAM_5K \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_5(10)  (.WCLK(\clk_2~O ), 
            .WE(\edb_top/la0/la_biu_inst/fifo_with_read_inst/we ), .WCLKE(1'b1), 
            .RCLK(\clk_2~O ), .RE(\edb_top/la0/la_biu_inst/fifo_with_read_inst/n136 ), 
            .WDATA({\edb_top/la0/cap_fifo_din_tu[4]_2 , \edb_top/la0/cap_fifo_din_tu[3]_2 , 
            \edb_top/la0/cap_fifo_din_tu[2]_2 , \edb_top/la0/cap_fifo_din_tu[1]_2 , 
            \edb_top/la0/cap_fifo_din_tu[0]_2 }), .WADDR({\edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]_2 , 
            \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]_2 , 
            \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]_2 , 
            \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]_2 , 
            \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]_2 , 
            \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]_2 , 
            \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]_2 , 
            \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]_2 , 
            \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]_2 , 
            \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]_2 }), 
            .RADDR({\edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , \edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , \edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , \edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , \edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), .RDATA({\edb_top/la0/la_biu_inst/swapped_data_out[4] , 
            \edb_top/la0/la_biu_inst/swapped_data_out[3] , \edb_top/la0/la_biu_inst/swapped_data_out[2] , 
            \edb_top/la0/la_biu_inst/swapped_data_out[1] , \edb_top/la0/la_biu_inst/swapped_data_out[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(399)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_5(10) .READ_WIDTH = 5;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_5(10) .WRITE_WIDTH = 5;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_5(10) .WCLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_5(10) .WCLKE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_5(10) .WE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_5(10) .RCLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_5(10) .RE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_5(10) .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_5(10) .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_5(10) .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_5(10) .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_5(10) .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_5(10) .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_5(10) .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_5(10) .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_5(10) .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_5(10) .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_5(10) .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_5(10) .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_5(10) .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_5(10) .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_5(10) .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_5(10) .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_5(10) .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_5(10) .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_5(10) .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_5(10) .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_5(10) .OUTPUT_REG = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_5(10) .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_3(01)  (.WCLK(\clk_2~O ), 
            .WE(\edb_top/la0/la_biu_inst/fifo_with_read_inst/we ), .WCLKE(1'b1), 
            .RCLK(\clk_2~O ), .RE(\edb_top/la0/la_biu_inst/fifo_with_read_inst/n136 ), 
            .WDATA({Open_0, \edb_top/la0/cap_fifo_din_tu[7]_2 , \edb_top/la0/cap_fifo_din_tu[6]_2 , 
            \edb_top/la0/cap_fifo_din_tu[5]_2 }), .WADDR({\edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]_2 , 
            \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]_2 , 
            \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]_2 , 
            \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]_2 , 
            \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]_2 , 
            \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]_2 , 
            \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]_2 , 
            \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]_2 , 
            \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]_2 , 
            \edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]_2 }), 
            .RADDR({\edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , \edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , \edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , \edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , \edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), .RDATA({Open_1, 
            \edb_top/la0/la_biu_inst/swapped_data_out[7] , \edb_top/la0/la_biu_inst/swapped_data_out[6] , 
            \edb_top/la0/la_biu_inst/swapped_data_out[5] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=4, WRITE_WIDTH=4, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000 */ ;   // C:/Efinity/2019.3/project/demo_led_loop/FPGA_prj/led_loop/debug_top.v(399)
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_3(01) .READ_WIDTH = 4;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_3(01) .WRITE_WIDTH = 4;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_3(01) .WCLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_3(01) .WCLKE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_3(01) .WE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_3(01) .RCLK_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_3(01) .RE_POLARITY = 1'b1;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_3(01) .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_3(01) .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_3(01) .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_3(01) .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_3(01) .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_3(01) .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_3(01) .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_3(01) .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_3(01) .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_3(01) .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_3(01) .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_3(01) .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_3(01) .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_3(01) .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_3(01) .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_3(01) .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_3(01) .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_3(01) .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_3(01) .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_3(01) .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_3(01) .OUTPUT_REG = 1'b0;
    defparam \edb_top/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__10_3(01) .WRITE_MODE = "READ_FIRST";
    EFX_LUT4 LUT__2646 (.I0(\edb_top/la0/module_state[2] ), .I1(\edb_top/la0/module_state[3] ), 
            .I2(\edb_top/la0/module_state[1] ), .O(n1685)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__2646.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__2647 (.I0(\edb_top/la0/module_state[3] ), .I1(\edb_top/la0/biu_ready ), 
            .I2(bscan_UPDATE), .I3(\edb_top/la0/module_state[1] ), .O(n1686)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__2647.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__2648 (.I0(n1684), .I1(n1686), .I2(\edb_top/la0/module_state[0] ), 
            .I3(n1685), .O(n1687)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__2648.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__2649 (.I0(\edb_top/la0/module_state[0] ), .I1(\edb_top/la0/module_state[1] ), 
            .I2(\edb_top/la0/module_state[2] ), .I3(\edb_top/la0/module_state[3] ), 
            .O(n1688)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__2649.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__2650 (.I0(\edb_top/edb_user_dr[81] ), .I1(n1688), .I2(bscan_UPDATE), 
            .I3(n1683), .O(n1689)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__2650.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__2651 (.I0(\edb_top/edb_user_dr[77] ), .I1(\edb_top/edb_user_dr[78] ), 
            .I2(\edb_top/edb_user_dr[79] ), .I3(\edb_top/edb_user_dr[80] ), 
            .O(n1690)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe1f */ ;
    defparam LUT__2651.LUTMASK = 16'hfe1f;
    EFX_LUT4 LUT__2652 (.I0(n1690), .I1(n1689), .O(n990)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__2652.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__2653 (.I0(\edb_top/la0/bit_count[0] ), .I1(\edb_top/la0/bit_count[1] ), 
            .I2(\edb_top/la0/bit_count[2] ), .O(n1691)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__2653.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__2654 (.I0(\edb_top/la0/bit_count[3] ), .I1(\edb_top/la0/bit_count[4] ), 
            .I2(n1691), .I3(\edb_top/la0/bit_count[5] ), .O(n1692)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__2654.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__2655 (.I0(\edb_top/la0/word_count[11] ), .I1(\edb_top/la0/word_count[12] ), 
            .I2(\edb_top/la0/word_count[13] ), .I3(\edb_top/la0/word_count[14] ), 
            .O(n1693)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__2655.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__2656 (.I0(\edb_top/la0/word_count[8] ), .I1(\edb_top/la0/word_count[9] ), 
            .I2(\edb_top/la0/word_count[10] ), .I3(\edb_top/la0/word_count[15] ), 
            .O(n1694)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__2656.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__2657 (.I0(\edb_top/la0/word_count[3] ), .I1(\edb_top/la0/word_count[4] ), 
            .I2(\edb_top/la0/word_count[5] ), .I3(\edb_top/la0/word_count[6] ), 
            .O(n1695)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__2657.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__2658 (.I0(\edb_top/la0/word_count[0] ), .I1(\edb_top/la0/word_count[1] ), 
            .I2(\edb_top/la0/word_count[2] ), .I3(\edb_top/la0/word_count[7] ), 
            .O(n1696)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__2658.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__2659 (.I0(n1693), .I1(n1694), .I2(n1695), .I3(n1696), 
            .O(n1697)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2659.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2660 (.I0(n1692), .I1(n1697), .I2(\edb_top/la0/module_state[0] ), 
            .I3(\edb_top/la0/module_state[1] ), .O(n1698)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h050c */ ;
    defparam LUT__2660.LUTMASK = 16'h050c;
    EFX_LUT4 LUT__2661 (.I0(\edb_top/la0/module_state[2] ), .I1(\edb_top/la0/module_state[3] ), 
            .O(n1699)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__2661.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__2662 (.I0(bscan_UPDATE), .I1(n1699), .O(n1700)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__2662.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__2663 (.I0(n1698), .I1(n1700), .I2(n1687), .I3(n990), 
            .O(n1701)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__2663.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__2664 (.I0(\edb_top/la0/module_state[0] ), .I1(\edb_top/la0/module_state[1] ), 
            .I2(n1701), .I3(n1699), .O(n1702)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf00 */ ;
    defparam LUT__2664.LUTMASK = 16'hbf00;
    EFX_LUT4 LUT__2665 (.I0(\edb_top/la0/crc_data_out[17] ), .I1(\edb_top/edb_user_dr[67] ), 
            .I2(\edb_top/la0/crc_data_out[23] ), .I3(\edb_top/edb_user_dr[73] ), 
            .O(n1703)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__2665.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__2666 (.I0(\edb_top/la0/crc_data_out[2] ), .I1(\edb_top/edb_user_dr[52] ), 
            .I2(\edb_top/la0/crc_data_out[28] ), .I3(\edb_top/edb_user_dr[78] ), 
            .O(n1704)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__2666.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__2667 (.I0(\edb_top/la0/crc_data_out[7] ), .I1(\edb_top/edb_user_dr[57] ), 
            .I2(\edb_top/la0/crc_data_out[31] ), .I3(\edb_top/edb_user_dr[81] ), 
            .O(n1705)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__2667.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__2668 (.I0(\edb_top/la0/crc_data_out[4] ), .I1(\edb_top/edb_user_dr[54] ), 
            .I2(\edb_top/la0/crc_data_out[21] ), .I3(\edb_top/edb_user_dr[71] ), 
            .O(n1706)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__2668.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__2669 (.I0(n1703), .I1(n1704), .I2(n1705), .I3(n1706), 
            .O(n1707)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2669.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2670 (.I0(\edb_top/la0/crc_data_out[8] ), .I1(\edb_top/edb_user_dr[58] ), 
            .I2(\edb_top/la0/crc_data_out[25] ), .I3(\edb_top/edb_user_dr[75] ), 
            .O(n1708)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__2670.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__2671 (.I0(\edb_top/la0/crc_data_out[10] ), .I1(\edb_top/edb_user_dr[60] ), 
            .I2(\edb_top/la0/crc_data_out[27] ), .I3(\edb_top/edb_user_dr[77] ), 
            .O(n1709)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__2671.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__2672 (.I0(\edb_top/la0/crc_data_out[12] ), .I1(\edb_top/edb_user_dr[62] ), 
            .I2(\edb_top/la0/crc_data_out[15] ), .I3(\edb_top/edb_user_dr[65] ), 
            .O(n1710)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__2672.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__2673 (.I0(\edb_top/la0/crc_data_out[18] ), .I1(\edb_top/edb_user_dr[68] ), 
            .I2(\edb_top/la0/crc_data_out[26] ), .I3(\edb_top/edb_user_dr[76] ), 
            .O(n1711)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__2673.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__2674 (.I0(n1708), .I1(n1709), .I2(n1710), .I3(n1711), 
            .O(n1712)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2674.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2675 (.I0(\edb_top/la0/crc_data_out[6] ), .I1(\edb_top/edb_user_dr[56] ), 
            .I2(\edb_top/la0/crc_data_out[11] ), .I3(\edb_top/edb_user_dr[61] ), 
            .O(n1713)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__2675.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__2676 (.I0(\edb_top/la0/crc_data_out[13] ), .I1(\edb_top/edb_user_dr[63] ), 
            .I2(\edb_top/la0/crc_data_out[19] ), .I3(\edb_top/edb_user_dr[69] ), 
            .O(n1714)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__2676.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__2677 (.I0(\edb_top/la0/crc_data_out[16] ), .I1(\edb_top/edb_user_dr[66] ), 
            .I2(\edb_top/la0/crc_data_out[24] ), .I3(\edb_top/edb_user_dr[74] ), 
            .O(n1715)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__2677.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__2678 (.I0(\edb_top/la0/crc_data_out[3] ), .I1(\edb_top/edb_user_dr[53] ), 
            .I2(\edb_top/la0/crc_data_out[29] ), .I3(\edb_top/edb_user_dr[79] ), 
            .O(n1716)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__2678.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__2679 (.I0(n1713), .I1(n1714), .I2(n1715), .I3(n1716), 
            .O(n1717)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2679.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2680 (.I0(\edb_top/la0/crc_data_out[0] ), .I1(\edb_top/edb_user_dr[50] ), 
            .I2(\edb_top/la0/crc_data_out[9] ), .I3(\edb_top/edb_user_dr[59] ), 
            .O(n1718)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__2680.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__2681 (.I0(\edb_top/la0/crc_data_out[5] ), .I1(\edb_top/edb_user_dr[55] ), 
            .I2(\edb_top/la0/crc_data_out[14] ), .I3(\edb_top/edb_user_dr[64] ), 
            .O(n1719)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__2681.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__2682 (.I0(\edb_top/la0/crc_data_out[20] ), .I1(\edb_top/edb_user_dr[70] ), 
            .I2(\edb_top/la0/crc_data_out[30] ), .I3(\edb_top/edb_user_dr[80] ), 
            .O(n1720)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__2682.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__2683 (.I0(\edb_top/la0/crc_data_out[1] ), .I1(\edb_top/edb_user_dr[51] ), 
            .I2(\edb_top/la0/crc_data_out[22] ), .I3(\edb_top/edb_user_dr[72] ), 
            .O(n1721)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__2683.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__2684 (.I0(n1718), .I1(n1719), .I2(n1720), .I3(n1721), 
            .O(n1722)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2684.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2685 (.I0(n1707), .I1(n1712), .I2(n1717), .I3(n1722), 
            .O(n1723)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2685.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2686 (.I0(\edb_top/la0/crc_data_out[0] ), .I1(\edb_top/la0/module_state[0] ), 
            .I2(n1723), .I3(\edb_top/la0/module_state[1] ), .O(n1724)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0bb */ ;
    defparam LUT__2686.LUTMASK = 16'hf0bb;
    EFX_LUT4 LUT__2687 (.I0(\edb_top/la0/biu_ready ), .I1(\edb_top/la0/module_state[1] ), 
            .I2(\edb_top/la0/data_out_shift_reg[0] ), .I3(n1699), .O(n1725)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__2687.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__2688 (.I0(n532), .I1(n534), .I2(n574), .I3(n575), 
            .O(n1726)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__2688.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__2689 (.I0(n1725), .I1(\edb_top/la0/module_state[0] ), 
            .I2(n1726), .O(n1727)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__2689.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__2690 (.I0(\edb_top/la0/biu_ready ), .I1(\edb_top/la0/module_state[0] ), 
            .I2(\edb_top/la0/data_out_shift_reg[0] ), .I3(n1685), .O(n1728)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0 */ ;
    defparam LUT__2690.LUTMASK = 16'hbbf0;
    EFX_LUT4 LUT__2691 (.I0(n1724), .I1(n1728), .I2(n1702), .I3(n1727), 
            .O(bscan_TDO)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__2691.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__2692 (.I0(\cnt[22] ), .I1(\cnt[20] ), .I2(\cnt[21] ), 
            .I3(\cnt[19] ), .O(n1729)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__2692.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__2693 (.I0(\cnt[16] ), .I1(n1729), .I2(\cnt[17] ), .I3(\cnt[18] ), 
            .O(n1730)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__2693.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__2694 (.I0(\cnt[0] ), .I1(\cnt[1] ), .I2(\cnt[2] ), .I3(\cnt[30] ), 
            .O(n1731)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__2694.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__2695 (.I0(\cnt[3] ), .I1(\cnt[4] ), .I2(\cnt[6] ), .I3(\cnt[5] ), 
            .O(n1732)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__2695.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__2696 (.I0(\cnt[8] ), .I1(\cnt[9] ), .I2(\cnt[14] ), 
            .I3(\cnt[10] ), .O(n1733)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__2696.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__2697 (.I0(\cnt[7] ), .I1(\cnt[11] ), .I2(\cnt[12] ), 
            .I3(\cnt[13] ), .O(n1734)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__2697.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__2698 (.I0(n1731), .I1(n1732), .I2(n1733), .I3(n1734), 
            .O(n1735)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2698.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2699 (.I0(\cnt[24] ), .I1(\cnt[25] ), .I2(\cnt[26] ), 
            .I3(\cnt[15] ), .O(n1736)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__2699.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__2700 (.I0(\cnt[27] ), .I1(\cnt[28] ), .I2(\cnt[29] ), 
            .I3(\cnt[23] ), .O(n1737)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__2700.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__2701 (.I0(n1730), .I1(n1735), .I2(n1736), .I3(n1737), 
            .O(n969)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff */ ;
    defparam LUT__2701.LUTMASK = 16'h7fff;
    EFX_LUT4 LUT__2702 (.I0(n969), .I1(lock), .O(n972)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7777 */ ;
    defparam LUT__2702.LUTMASK = 16'h7777;
    EFX_LUT4 LUT__2703 (.I0(\edb_top/la0/module_state[1] ), .I1(\edb_top/la0/module_state[0] ), 
            .O(n1738)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__2703.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__2704 (.I0(n1699), .I1(n1738), .O(n1277)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2704.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2705 (.I0(n1277), .I1(\edb_top/edb_user_dr[42] ), .O(n973)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__2705.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__2706 (.I0(\edb_top/edb_user_dr[78] ), .I1(\edb_top/edb_user_dr[77] ), 
            .I2(n1689), .I3(\edb_top/edb_user_dr[80] ), .O(n1008)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__2706.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__2707 (.I0(\edb_top/edb_user_dr[71] ), .I1(\edb_top/edb_user_dr[75] ), 
            .I2(\edb_top/edb_user_dr[76] ), .I3(\edb_top/edb_user_dr[79] ), 
            .O(n1739)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__2707.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__2708 (.I0(\edb_top/edb_user_dr[72] ), .I1(\edb_top/edb_user_dr[73] ), 
            .I2(\edb_top/edb_user_dr[74] ), .I3(n1739), .O(n1740)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__2708.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__2709 (.I0(n1008), .I1(n1740), .O(n1741)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2709.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2710 (.I0(\edb_top/edb_user_dr[70] ), .I1(n1741), .O(n1742)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__2710.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__2711 (.I0(\edb_top/edb_user_dr[66] ), .I1(\edb_top/edb_user_dr[67] ), 
            .I2(\edb_top/edb_user_dr[68] ), .I3(\edb_top/edb_user_dr[69] ), 
            .O(n1743)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__2711.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__2712 (.I0(\edb_top/edb_user_dr[64] ), .I1(\edb_top/edb_user_dr[65] ), 
            .I2(n1743), .O(n1744)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__2712.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__2713 (.I0(n1742), .I1(n1744), .I2(n1277), .O(n975)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__2713.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__2714 (.I0(n1742), .I1(n1744), .O(n978)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2714.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2715 (.I0(n1277), .I1(\edb_top/edb_user_dr[43] ), .O(n979)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__2715.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__2716 (.I0(n1277), .I1(\edb_top/edb_user_dr[44] ), .O(n980)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__2716.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__2717 (.I0(\edb_top/edb_user_dr[65] ), .I1(n1743), .I2(\edb_top/edb_user_dr[64] ), 
            .I3(n1742), .O(n982)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__2717.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__2718 (.I0(\edb_top/la0/address_counter[7] ), .I1(\edb_top/la0/address_counter[8] ), 
            .I2(\edb_top/la0/address_counter[9] ), .I3(\edb_top/la0/address_counter[10] ), 
            .O(n1745)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__2718.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__2719 (.I0(\edb_top/la0/address_counter[11] ), .I1(\edb_top/la0/address_counter[12] ), 
            .I2(\edb_top/la0/address_counter[13] ), .I3(n1745), .O(n1746)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__2719.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__2720 (.I0(\edb_top/la0/address_counter[3] ), .I1(\edb_top/la0/address_counter[4] ), 
            .I2(\edb_top/la0/address_counter[5] ), .I3(\edb_top/la0/address_counter[14] ), 
            .O(n1747)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__2720.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__2721 (.I0(\edb_top/la0/address_counter[0] ), .I1(\edb_top/la0/address_counter[1] ), 
            .I2(\edb_top/la0/address_counter[2] ), .I3(\edb_top/la0/address_counter[6] ), 
            .O(n1748)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__2721.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__2722 (.I0(n1746), .I1(n1747), .I2(n1748), .O(n1749)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__2722.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__2723 (.I0(n1749), .I1(n34), .I2(\edb_top/edb_user_dr[45] ), 
            .I3(n1688), .O(n983)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044 */ ;
    defparam LUT__2723.LUTMASK = 16'hf044;
    EFX_LUT4 LUT__2724 (.I0(\edb_top/la0/opcode[1] ), .I1(\edb_top/la0/opcode[3] ), 
            .I2(\edb_top/la0/opcode[2] ), .I3(\edb_top/la0/opcode[0] ), 
            .O(n986)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__2724.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__2725 (.I0(\edb_top/la0/bit_count[0] ), .I1(\edb_top/la0/bit_count[1] ), 
            .I2(\edb_top/la0/bit_count[2] ), .O(n1750)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__2725.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__2726 (.I0(\edb_top/la0/bit_count[3] ), .I1(\edb_top/la0/bit_count[4] ), 
            .I2(\edb_top/la0/bit_count[5] ), .O(n1751)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__2726.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__2727 (.I0(n1691), .I1(n1750), .I2(n986), .I3(n1751), 
            .O(n1752)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__2727.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__2728 (.I0(\edb_top/la0/module_state[3] ), .I1(\edb_top/la0/module_state[2] ), 
            .O(n1753)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__2728.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__2729 (.I0(\edb_top/la0/module_state[0] ), .I1(\edb_top/la0/module_state[1] ), 
            .I2(n1752), .I3(n1753), .O(n1754)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__2729.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__2730 (.I0(n678), .I1(n680), .I2(n682), .I3(n684), 
            .O(n1755)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__2730.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__2731 (.I0(n672), .I1(n674), .I2(n676), .I3(n686), 
            .O(n1756)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__2731.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__2732 (.I0(n662), .I1(n664), .I2(n666), .I3(n668), 
            .O(n1757)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__2732.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__2733 (.I0(n40), .I1(n659), .I2(n660), .I3(n670), .O(n1758)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__2733.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__2734 (.I0(n1755), .I1(n1756), .I2(n1757), .I3(n1758), 
            .O(n1759)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2734.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2735 (.I0(n1697), .I1(n1759), .I2(\edb_top/la0/module_state[0] ), 
            .O(n1760)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__2735.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__2736 (.I0(n1760), .I1(n1754), .I2(\edb_top/la0/module_state[2] ), 
            .I3(\edb_top/la0/module_state[3] ), .O(n1761)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbb0 */ ;
    defparam LUT__2736.LUTMASK = 16'hbbb0;
    EFX_LUT4 LUT__2737 (.I0(bscan_UPDATE), .I1(n1685), .I2(\edb_top/la0/module_state[0] ), 
            .I3(\edb_top/la0/biu_ready ), .O(n1762)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__2737.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__2738 (.I0(n1759), .I1(n1762), .I2(n1738), .O(n1763)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__2738.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__2739 (.I0(n1763), .I1(n1697), .I2(\edb_top/la0/module_state[2] ), 
            .O(n1764)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__2739.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__2740 (.I0(\edb_top/la0/module_state[0] ), .I1(\edb_top/la0/module_state[1] ), 
            .O(n1765)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__2740.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__2741 (.I0(n1765), .I1(n1764), .I2(n1761), .O(n1766)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7c7c */ ;
    defparam LUT__2741.LUTMASK = 16'h7c7c;
    EFX_LUT4 LUT__2742 (.I0(n990), .I1(n1766), .O(n984)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__2742.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__2743 (.I0(n990), .I1(n1699), .O(n1767)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__2743.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__2744 (.I0(n1767), .I1(n1765), .I2(n1762), .I3(n1754), 
            .O(n1768)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__2744.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__2745 (.I0(\edb_top/la0/bit_count[0] ), .I1(n1768), .O(n991)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__2745.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__2746 (.I0(bscan_UPDATE), .I1(\edb_top/la0/module_state[0] ), 
            .O(n1769)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__2746.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__2747 (.I0(n1683), .I1(\edb_top/edb_user_dr[81] ), .I2(n1769), 
            .I3(\edb_top/la0/module_state[1] ), .O(n1770)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00 */ ;
    defparam LUT__2747.LUTMASK = 16'h7f00;
    EFX_LUT4 LUT__2748 (.I0(n1770), .I1(\edb_top/la0/module_state[0] ), 
            .I2(n1753), .O(n1771)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090 */ ;
    defparam LUT__2748.LUTMASK = 16'h9090;
    EFX_LUT4 LUT__2749 (.I0(n1767), .I1(\edb_top/la0/module_state[0] ), 
            .I2(n1762), .I3(n1771), .O(n992)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e */ ;
    defparam LUT__2749.LUTMASK = 16'h000e;
    EFX_LUT4 LUT__2750 (.I0(\edb_top/edb_user_dr[29] ), .I1(n40), .I2(n1688), 
            .O(n994)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__2750.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__2751 (.I0(n1697), .I1(n1752), .O(n1772)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2751.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2752 (.I0(n1684), .I1(n1697), .I2(\edb_top/la0/module_state[0] ), 
            .I3(\edb_top/la0/module_state[1] ), .O(n1773)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__2752.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__2753 (.I0(n1769), .I1(n1772), .I2(n1773), .I3(n1753), 
            .O(n1774)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__2753.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__2754 (.I0(\edb_top/la0/module_state[0] ), .I1(n1770), 
            .I2(n1774), .I3(n1768), .O(n995)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h10ff */ ;
    defparam LUT__2754.LUTMASK = 16'h10ff;
    EFX_LUT4 LUT__2755 (.I0(\edb_top/la0/internal_register_select[2] ), .I1(\edb_top/la0/internal_register_select[3] ), 
            .I2(\edb_top/la0/internal_register_select[4] ), .I3(\edb_top/la0/internal_register_select[5] ), 
            .O(n1775)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__2755.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__2756 (.I0(\edb_top/la0/internal_register_select[0] ), .I1(\edb_top/la0/internal_register_select[1] ), 
            .I2(n1775), .I3(\edb_top/la0/internal_register_select[6] ), 
            .O(n1776)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__2756.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__2757 (.I0(\edb_top/la0/internal_register_select[0] ), .I1(n1775), 
            .I2(\edb_top/la0/internal_register_select[1] ), .I3(\edb_top/la0/internal_register_select[6] ), 
            .O(n1777)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__2757.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__2758 (.I0(n1776), .I1(\edb_top/la0/register_conn[64][0] ), 
            .I2(n1777), .I3(\edb_top/la0/register_conn[66][0] ), .O(n1778)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2758.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2759 (.I0(\edb_top/la0/internal_register_select[0] ), .I1(\edb_top/la0/internal_register_select[1] ), 
            .I2(\edb_top/la0/internal_register_select[6] ), .I3(n1775), 
            .O(n1779)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__2759.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__2760 (.I0(n1779), .I1(\edb_top/la0/register_conn[0][0] ), 
            .I2(n1778), .O(n1780)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2760.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2761 (.I0(bscan_UPDATE), .I1(\edb_top/la0/module_state[0] ), 
            .I2(\edb_top/la0/module_state[1] ), .I3(\edb_top/la0/biu_ready ), 
            .O(n1781)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__2761.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__2762 (.I0(n1781), .I1(n1765), .I2(\edb_top/la0/module_state[2] ), 
            .O(n1782)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3d3d */ ;
    defparam LUT__2762.LUTMASK = 16'h3d3d;
    EFX_LUT4 LUT__2763 (.I0(\edb_top/la0/internal_register_select[8] ), .I1(\edb_top/la0/internal_register_select[9] ), 
            .I2(\edb_top/la0/internal_register_select[10] ), .I3(\edb_top/la0/internal_register_select[11] ), 
            .O(n1783)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__2763.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__2764 (.I0(\edb_top/la0/internal_register_select[7] ), .I1(\edb_top/la0/internal_register_select[12] ), 
            .I2(n1783), .O(n1784)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__2764.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__2765 (.I0(n1782), .I1(n1784), .O(n1785)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2765.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2766 (.I0(\edb_top/la0/internal_register_select[1] ), .I1(\edb_top/la0/internal_register_select[6] ), 
            .I2(n1775), .I3(\edb_top/la0/internal_register_select[0] ), 
            .O(n1786)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__2766.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__2767 (.I0(\edb_top/la0/la_trig_mask[0] ), .I1(n1786), 
            .I2(n1780), .I3(n1785), .O(n1787)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__2767.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__2768 (.I0(n1752), .I1(\edb_top/la0/module_state[2] ), 
            .O(n1788)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__2768.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__2769 (.I0(n1683), .I1(n1765), .I2(bscan_CAPTURE), .O(n1789)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__2769.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__2770 (.I0(n1782), .I1(n1789), .I2(n1788), .I3(\edb_top/la0/module_state[3] ), 
            .O(n1790)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__2770.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__2771 (.I0(\edb_top/la0/module_state[3] ), .I1(n1784), 
            .I2(n1789), .I3(n1782), .O(n1791)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__2771.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__2772 (.I0(\edb_top/la0/internal_register_select[1] ), .I1(\edb_top/la0/internal_register_select[0] ), 
            .I2(n1775), .I3(\edb_top/la0/internal_register_select[6] ), 
            .O(n1792)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__2772.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__2773 (.I0(n1791), .I1(n1792), .I2(\edb_top/la0/register_conn[65][0] ), 
            .O(n1793)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__2773.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__2774 (.I0(n1782), .I1(\edb_top/la0/data_from_biu[0] ), 
            .I2(n1790), .I3(n1793), .O(n1794)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf */ ;
    defparam LUT__2774.LUTMASK = 16'h00bf;
    EFX_LUT4 LUT__2775 (.I0(n1787), .I1(\edb_top/la0/data_out_shift_reg[1] ), 
            .I2(n1790), .I3(n1794), .O(n996)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacff */ ;
    defparam LUT__2775.LUTMASK = 16'hacff;
    EFX_LUT4 LUT__2776 (.I0(n1683), .I1(bscan_SHIFT), .I2(\edb_top/la0/module_state[2] ), 
            .O(n1795)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__2776.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__2777 (.I0(\edb_top/la0/module_state[3] ), .I1(n1795), 
            .I2(n1765), .I3(n1790), .O(n997)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__2777.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__2778 (.I0(bscan_UPDATE), .I1(n1772), .I2(\edb_top/la0/module_state[0] ), 
            .I3(n1770), .O(n1796)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__2778.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__2779 (.I0(n1796), .I1(n1774), .I2(n1701), .O(n998)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f4f */ ;
    defparam LUT__2779.LUTMASK = 16'h4f4f;
    EFX_LUT4 LUT__2780 (.I0(n1741), .I1(\edb_top/edb_user_dr[70] ), .O(n1797)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2780.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2781 (.I0(n1797), .I1(n1744), .O(n1001)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2781.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2782 (.I0(\edb_top/edb_user_dr[65] ), .I1(n1743), .I2(\edb_top/edb_user_dr[64] ), 
            .I3(n1797), .O(n1002)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__2782.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__2783 (.I0(\edb_top/edb_user_dr[64] ), .I1(n1743), .I2(n1797), 
            .I3(\edb_top/edb_user_dr[65] ), .O(n1003)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__2783.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__2784 (.I0(n1749), .I1(n756), .I2(\edb_top/edb_user_dr[46] ), 
            .I3(n1688), .O(n1071)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044 */ ;
    defparam LUT__2784.LUTMASK = 16'hf044;
    EFX_LUT4 LUT__2785 (.I0(n1749), .I1(n754), .I2(\edb_top/edb_user_dr[47] ), 
            .I3(n1688), .O(n1072)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044 */ ;
    defparam LUT__2785.LUTMASK = 16'hf044;
    EFX_LUT4 LUT__2786 (.I0(n1749), .I1(n752), .I2(\edb_top/edb_user_dr[48] ), 
            .I3(n1688), .O(n1073)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044 */ ;
    defparam LUT__2786.LUTMASK = 16'hf044;
    EFX_LUT4 LUT__2787 (.I0(n1749), .I1(n750), .I2(\edb_top/edb_user_dr[49] ), 
            .I3(n1688), .O(n1074)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044 */ ;
    defparam LUT__2787.LUTMASK = 16'hf044;
    EFX_LUT4 LUT__2788 (.I0(n1749), .I1(n748), .I2(\edb_top/edb_user_dr[50] ), 
            .I3(n1688), .O(n1075)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044 */ ;
    defparam LUT__2788.LUTMASK = 16'hf044;
    EFX_LUT4 LUT__2789 (.I0(n1749), .I1(n746), .I2(\edb_top/edb_user_dr[51] ), 
            .I3(n1688), .O(n1076)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044 */ ;
    defparam LUT__2789.LUTMASK = 16'hf044;
    EFX_LUT4 LUT__2790 (.I0(n1749), .I1(n744), .I2(\edb_top/edb_user_dr[52] ), 
            .I3(n1688), .O(n1077)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044 */ ;
    defparam LUT__2790.LUTMASK = 16'hf044;
    EFX_LUT4 LUT__2791 (.I0(n1749), .I1(n742), .I2(\edb_top/edb_user_dr[53] ), 
            .I3(n1688), .O(n1078)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044 */ ;
    defparam LUT__2791.LUTMASK = 16'hf044;
    EFX_LUT4 LUT__2792 (.I0(n1749), .I1(n740), .I2(\edb_top/edb_user_dr[54] ), 
            .I3(n1688), .O(n1079)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044 */ ;
    defparam LUT__2792.LUTMASK = 16'hf044;
    EFX_LUT4 LUT__2793 (.I0(n1749), .I1(n738), .I2(\edb_top/edb_user_dr[55] ), 
            .I3(n1688), .O(n1080)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044 */ ;
    defparam LUT__2793.LUTMASK = 16'hf044;
    EFX_LUT4 LUT__2794 (.I0(n1749), .I1(n736), .I2(\edb_top/edb_user_dr[56] ), 
            .I3(n1688), .O(n1081)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044 */ ;
    defparam LUT__2794.LUTMASK = 16'hf044;
    EFX_LUT4 LUT__2795 (.I0(n1749), .I1(n734), .I2(\edb_top/edb_user_dr[57] ), 
            .I3(n1688), .O(n1082)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044 */ ;
    defparam LUT__2795.LUTMASK = 16'hf044;
    EFX_LUT4 LUT__2796 (.I0(n1749), .I1(n732), .I2(\edb_top/edb_user_dr[58] ), 
            .I3(n1688), .O(n1083)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044 */ ;
    defparam LUT__2796.LUTMASK = 16'hf044;
    EFX_LUT4 LUT__2797 (.I0(n1749), .I1(n730), .I2(\edb_top/edb_user_dr[59] ), 
            .I3(n1688), .O(n1084)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044 */ ;
    defparam LUT__2797.LUTMASK = 16'hf044;
    EFX_LUT4 LUT__2798 (.I0(\edb_top/la0/address_counter[15] ), .I1(n728), 
            .I2(n1749), .O(n1798)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__2798.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__2799 (.I0(n1798), .I1(\edb_top/edb_user_dr[60] ), .I2(n1688), 
            .O(n1085)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__2799.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__2800 (.I0(n24), .I1(n726), .I2(n1749), .O(n1799)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__2800.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__2801 (.I0(n1799), .I1(\edb_top/edb_user_dr[61] ), .I2(n1688), 
            .O(n1086)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__2801.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__2802 (.I0(n785), .I1(n724), .I2(n1749), .O(n1800)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__2802.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__2803 (.I0(n1800), .I1(\edb_top/edb_user_dr[62] ), .I2(n1688), 
            .O(n1087)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__2803.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__2804 (.I0(n783), .I1(n722), .I2(n1749), .O(n1801)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__2804.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__2805 (.I0(n1801), .I1(\edb_top/edb_user_dr[63] ), .I2(n1688), 
            .O(n1088)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__2805.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__2806 (.I0(n781), .I1(n720), .I2(n1749), .O(n1802)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__2806.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__2807 (.I0(n1802), .I1(\edb_top/edb_user_dr[64] ), .I2(n1688), 
            .O(n1089)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__2807.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__2808 (.I0(n779), .I1(n718), .I2(n1749), .O(n1803)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__2808.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__2809 (.I0(n1803), .I1(\edb_top/edb_user_dr[65] ), .I2(n1688), 
            .O(n1090)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__2809.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__2810 (.I0(n777), .I1(n716), .I2(n1749), .O(n1804)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__2810.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__2811 (.I0(n1804), .I1(\edb_top/edb_user_dr[66] ), .I2(n1688), 
            .O(n1091)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__2811.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__2812 (.I0(n775), .I1(n714), .I2(n1749), .O(n1805)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__2812.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__2813 (.I0(n1805), .I1(\edb_top/edb_user_dr[67] ), .I2(n1688), 
            .O(n1092)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__2813.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__2814 (.I0(n773), .I1(n712), .I2(n1749), .O(n1806)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__2814.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__2815 (.I0(n1806), .I1(\edb_top/edb_user_dr[68] ), .I2(n1688), 
            .O(n1093)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__2815.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__2816 (.I0(n771), .I1(n710), .I2(n1749), .O(n1807)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__2816.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__2817 (.I0(n1807), .I1(\edb_top/edb_user_dr[69] ), .I2(n1688), 
            .O(n1094)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__2817.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__2832 (.I0(n1768), .I1(n36), .O(n1105)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2832.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2833 (.I0(n1768), .I1(n695), .O(n1106)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2833.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2834 (.I0(n1768), .I1(n693), .O(n1107)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2834.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2835 (.I0(n1768), .I1(n691), .O(n1108)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2835.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2836 (.I0(n1768), .I1(n689), .O(n1109)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2836.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2837 (.I0(\edb_top/edb_user_dr[30] ), .I1(n686), .I2(n1688), 
            .O(n1110)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__2837.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__2838 (.I0(\edb_top/edb_user_dr[31] ), .I1(n684), .I2(n1688), 
            .O(n1111)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__2838.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__2839 (.I0(\edb_top/edb_user_dr[32] ), .I1(n682), .I2(n1688), 
            .O(n1112)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__2839.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__2840 (.I0(\edb_top/edb_user_dr[33] ), .I1(n680), .I2(n1688), 
            .O(n1113)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__2840.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__2841 (.I0(\edb_top/edb_user_dr[34] ), .I1(n678), .I2(n1688), 
            .O(n1114)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__2841.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__2842 (.I0(\edb_top/edb_user_dr[35] ), .I1(n676), .I2(n1688), 
            .O(n1115)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__2842.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__2843 (.I0(\edb_top/edb_user_dr[36] ), .I1(n674), .I2(n1688), 
            .O(n1116)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__2843.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__2844 (.I0(\edb_top/edb_user_dr[37] ), .I1(n672), .I2(n1688), 
            .O(n1117)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__2844.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__2845 (.I0(\edb_top/edb_user_dr[38] ), .I1(n670), .I2(n1688), 
            .O(n1118)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__2845.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__2846 (.I0(\edb_top/edb_user_dr[39] ), .I1(n668), .I2(n1688), 
            .O(n1119)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__2846.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__2847 (.I0(\edb_top/edb_user_dr[40] ), .I1(n666), .I2(n1688), 
            .O(n1120)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__2847.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__2848 (.I0(\edb_top/edb_user_dr[41] ), .I1(n664), .I2(n1688), 
            .O(n1121)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__2848.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__2849 (.I0(\edb_top/edb_user_dr[42] ), .I1(n662), .I2(n1688), 
            .O(n1122)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__2849.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__2850 (.I0(\edb_top/edb_user_dr[43] ), .I1(n660), .I2(n1688), 
            .O(n1123)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__2850.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__2851 (.I0(\edb_top/edb_user_dr[44] ), .I1(n659), .I2(n1688), 
            .O(n1124)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__2851.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__2852 (.I0(n1782), .I1(\edb_top/la0/data_from_biu[1] ), 
            .I2(\edb_top/la0/data_out_shift_reg[2] ), .I3(n1790), .O(n1815)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__2852.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__2853 (.I0(n1776), .I1(\edb_top/la0/register_conn[64][1] ), 
            .I2(n1777), .I3(\edb_top/la0/register_conn[66][1] ), .O(n1816)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2853.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2854 (.I0(n1786), .I1(\edb_top/la0/la_trig_mask[1] ), 
            .I2(n1792), .I3(\edb_top/la0/register_conn[65][1] ), .O(n1817)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2854.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2855 (.I0(n1779), .I1(\edb_top/la0/register_conn[0][1] ), 
            .I2(n1816), .I3(n1817), .O(n1818)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7000 */ ;
    defparam LUT__2855.LUTMASK = 16'h7000;
    EFX_LUT4 LUT__2856 (.I0(n1818), .I1(n1791), .I2(n1815), .O(n1125)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f4f */ ;
    defparam LUT__2856.LUTMASK = 16'h4f4f;
    EFX_LUT4 LUT__2857 (.I0(n1782), .I1(\edb_top/la0/data_from_biu[2] ), 
            .I2(\edb_top/la0/data_out_shift_reg[3] ), .I3(n1790), .O(n1819)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__2857.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__2858 (.I0(n1776), .I1(\edb_top/la0/register_conn[64][2] ), 
            .I2(n1777), .I3(\edb_top/la0/register_conn[66][2] ), .O(n1820)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2858.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2859 (.I0(n1786), .I1(\edb_top/la0/la_trig_mask[2] ), 
            .I2(n1792), .I3(\edb_top/la0/register_conn[65][2] ), .O(n1821)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2859.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2860 (.I0(n1779), .I1(\edb_top/la0/register_conn[0][2] ), 
            .I2(n1820), .I3(n1821), .O(n1822)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7000 */ ;
    defparam LUT__2860.LUTMASK = 16'h7000;
    EFX_LUT4 LUT__2861 (.I0(n1822), .I1(n1791), .I2(n1819), .O(n1126)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f4f */ ;
    defparam LUT__2861.LUTMASK = 16'h4f4f;
    EFX_LUT4 LUT__2862 (.I0(n1782), .I1(\edb_top/la0/data_from_biu[3] ), 
            .I2(\edb_top/la0/data_out_shift_reg[4] ), .I3(n1790), .O(n1823)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__2862.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__2863 (.I0(n1779), .I1(\edb_top/la0/la_run_trig ), .I2(n1777), 
            .I3(\edb_top/la0/register_conn[66][3] ), .O(n1824)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2863.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2864 (.I0(n1792), .I1(\edb_top/la0/register_conn[65][3] ), 
            .I2(n1824), .O(n1825)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2864.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2865 (.I0(n1786), .I1(\edb_top/la0/la_trig_mask[3] ), 
            .I2(n1825), .O(n1826)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2865.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2866 (.I0(n1826), .I1(n1791), .I2(n1823), .O(n1127)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f4f */ ;
    defparam LUT__2866.LUTMASK = 16'h4f4f;
    EFX_LUT4 LUT__2867 (.I0(n1782), .I1(\edb_top/la0/data_from_biu[4] ), 
            .I2(\edb_top/la0/data_out_shift_reg[5] ), .I3(n1790), .O(n1827)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__2867.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__2868 (.I0(n1779), .I1(\edb_top/la0/la_run_trig_imdt ), 
            .I2(n1777), .I3(\edb_top/la0/register_conn[66][4] ), .O(n1828)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2868.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2869 (.I0(n1792), .I1(\edb_top/la0/register_conn[65][4] ), 
            .I2(n1828), .O(n1829)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2869.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2870 (.I0(n1786), .I1(\edb_top/la0/la_trig_mask[4] ), 
            .I2(n1829), .O(n1830)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2870.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2871 (.I0(n1830), .I1(n1791), .I2(n1827), .O(n1128)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f4f */ ;
    defparam LUT__2871.LUTMASK = 16'h4f4f;
    EFX_LUT4 LUT__2872 (.I0(n1782), .I1(\edb_top/la0/data_from_biu[5] ), 
            .I2(\edb_top/la0/data_out_shift_reg[6] ), .I3(n1790), .O(n1831)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__2872.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__2873 (.I0(n1779), .I1(\edb_top/la0/la_stop_trig ), .I2(n1777), 
            .I3(\edb_top/la0/register_conn[66][5] ), .O(n1832)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2873.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2874 (.I0(n1792), .I1(\edb_top/la0/register_conn[65][5] ), 
            .I2(n1832), .O(n1833)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2874.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2875 (.I0(n1786), .I1(\edb_top/la0/la_trig_mask[5] ), 
            .I2(n1833), .O(n1834)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2875.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2876 (.I0(n1834), .I1(n1791), .I2(n1831), .O(n1129)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f4f */ ;
    defparam LUT__2876.LUTMASK = 16'h4f4f;
    EFX_LUT4 LUT__2877 (.I0(n1782), .I1(\edb_top/la0/data_from_biu[6] ), 
            .I2(\edb_top/la0/data_out_shift_reg[7] ), .I3(n1790), .O(n1835)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__2877.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__2878 (.I0(n1779), .I1(\edb_top/la0/la_trig_pos[0] ), .I2(n1777), 
            .I3(\edb_top/la0/register_conn[66][6] ), .O(n1836)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2878.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2879 (.I0(n1792), .I1(\edb_top/la0/register_conn[65][6] ), 
            .I2(n1836), .O(n1837)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2879.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2880 (.I0(n1786), .I1(\edb_top/la0/la_trig_mask[6] ), 
            .I2(n1837), .O(n1838)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2880.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2881 (.I0(n1838), .I1(n1791), .I2(n1835), .O(n1130)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f4f */ ;
    defparam LUT__2881.LUTMASK = 16'h4f4f;
    EFX_LUT4 LUT__2882 (.I0(n1782), .I1(\edb_top/la0/data_from_biu[7] ), 
            .I2(\edb_top/la0/data_out_shift_reg[8] ), .I3(n1790), .O(n1839)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__2882.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__2883 (.I0(n1779), .I1(\edb_top/la0/la_trig_pos[1] ), .I2(\edb_top/la0/register_conn[66][7] ), 
            .I3(n1777), .O(n1840)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2883.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2884 (.I0(n1792), .I1(\edb_top/la0/register_conn[65][7] ), 
            .I2(n1840), .O(n1841)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2884.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2885 (.I0(n1786), .I1(\edb_top/la0/la_trig_mask[7] ), 
            .I2(n1841), .O(n1842)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2885.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2886 (.I0(n1842), .I1(n1791), .I2(n1839), .O(n1131)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f4f */ ;
    defparam LUT__2886.LUTMASK = 16'h4f4f;
    EFX_LUT4 LUT__2887 (.I0(n1779), .I1(\edb_top/la0/la_trig_pos[2] ), .I2(\edb_top/la0/register_conn[66][8] ), 
            .I3(n1777), .O(n1843)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2887.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2888 (.I0(n1792), .I1(\edb_top/la0/register_conn[65][8] ), 
            .I2(n1843), .O(n1844)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2888.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2889 (.I0(n1786), .I1(\edb_top/la0/la_trig_mask[8] ), 
            .I2(n1844), .O(n1845)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2889.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2890 (.I0(n1845), .I1(n1791), .I2(n1790), .I3(\edb_top/la0/data_out_shift_reg[9] ), 
            .O(n1132)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44 */ ;
    defparam LUT__2890.LUTMASK = 16'h4f44;
    EFX_LUT4 LUT__2891 (.I0(n1779), .I1(\edb_top/la0/la_trig_pos[3] ), .I2(\edb_top/la0/register_conn[66][9] ), 
            .I3(n1777), .O(n1846)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2891.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2892 (.I0(n1792), .I1(\edb_top/la0/register_conn[65][9] ), 
            .I2(n1846), .O(n1847)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2892.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2893 (.I0(n1786), .I1(\edb_top/la0/la_trig_mask[9] ), 
            .I2(n1847), .O(n1848)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2893.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2894 (.I0(n1848), .I1(n1791), .I2(n1790), .I3(\edb_top/la0/data_out_shift_reg[10] ), 
            .O(n1133)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44 */ ;
    defparam LUT__2894.LUTMASK = 16'h4f44;
    EFX_LUT4 LUT__2895 (.I0(n1779), .I1(\edb_top/la0/la_trig_pos[4] ), .I2(\edb_top/la0/register_conn[66][10] ), 
            .I3(n1777), .O(n1849)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2895.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2896 (.I0(n1792), .I1(\edb_top/la0/register_conn[65][10] ), 
            .I2(n1849), .O(n1850)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2896.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2897 (.I0(n1786), .I1(\edb_top/la0/la_trig_mask[10] ), 
            .I2(n1850), .O(n1851)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2897.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2898 (.I0(n1851), .I1(n1791), .I2(n1790), .I3(\edb_top/la0/data_out_shift_reg[11] ), 
            .O(n1134)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44 */ ;
    defparam LUT__2898.LUTMASK = 16'h4f44;
    EFX_LUT4 LUT__2899 (.I0(n1779), .I1(\edb_top/la0/la_trig_pos[5] ), .I2(\edb_top/la0/register_conn[66][11] ), 
            .I3(n1777), .O(n1852)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2899.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2900 (.I0(n1792), .I1(\edb_top/la0/register_conn[65][11] ), 
            .I2(n1852), .O(n1853)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2900.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2901 (.I0(n1786), .I1(\edb_top/la0/la_trig_mask[11] ), 
            .I2(n1853), .O(n1854)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2901.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2902 (.I0(n1854), .I1(n1791), .I2(n1790), .I3(\edb_top/la0/data_out_shift_reg[12] ), 
            .O(n1135)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44 */ ;
    defparam LUT__2902.LUTMASK = 16'h4f44;
    EFX_LUT4 LUT__2903 (.I0(n1779), .I1(\edb_top/la0/la_trig_pos[6] ), .I2(\edb_top/la0/register_conn[66][12] ), 
            .I3(n1777), .O(n1855)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2903.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2904 (.I0(n1792), .I1(\edb_top/la0/register_conn[65][12] ), 
            .I2(n1855), .O(n1856)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2904.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2905 (.I0(n1786), .I1(\edb_top/la0/la_trig_mask[12] ), 
            .I2(n1856), .O(n1857)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2905.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2906 (.I0(n1857), .I1(n1791), .I2(n1790), .I3(\edb_top/la0/data_out_shift_reg[13] ), 
            .O(n1136)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44 */ ;
    defparam LUT__2906.LUTMASK = 16'h4f44;
    EFX_LUT4 LUT__2907 (.I0(n1779), .I1(\edb_top/la0/la_trig_pos[7] ), .I2(\edb_top/la0/register_conn[66][13] ), 
            .I3(n1777), .O(n1858)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2907.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2908 (.I0(n1792), .I1(\edb_top/la0/register_conn[65][13] ), 
            .I2(n1858), .O(n1859)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2908.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2909 (.I0(n1786), .I1(\edb_top/la0/la_trig_mask[13] ), 
            .I2(n1859), .O(n1860)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2909.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2910 (.I0(n1860), .I1(n1791), .I2(n1790), .I3(\edb_top/la0/data_out_shift_reg[14] ), 
            .O(n1137)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44 */ ;
    defparam LUT__2910.LUTMASK = 16'h4f44;
    EFX_LUT4 LUT__2911 (.I0(n1779), .I1(\edb_top/la0/la_trig_pos[8] ), .I2(\edb_top/la0/register_conn[66][14] ), 
            .I3(n1777), .O(n1861)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2911.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2912 (.I0(n1792), .I1(\edb_top/la0/register_conn[65][14] ), 
            .I2(n1861), .O(n1862)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2912.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2913 (.I0(n1786), .I1(\edb_top/la0/la_trig_mask[14] ), 
            .I2(n1862), .O(n1863)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2913.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2914 (.I0(n1863), .I1(n1791), .I2(n1790), .I3(\edb_top/la0/data_out_shift_reg[15] ), 
            .O(n1138)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44 */ ;
    defparam LUT__2914.LUTMASK = 16'h4f44;
    EFX_LUT4 LUT__2915 (.I0(n1779), .I1(\edb_top/la0/la_trig_pos[9] ), .I2(\edb_top/la0/register_conn[66][15] ), 
            .I3(n1777), .O(n1864)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2915.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2916 (.I0(n1792), .I1(\edb_top/la0/register_conn[65][15] ), 
            .I2(n1864), .O(n1865)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2916.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2917 (.I0(n1786), .I1(\edb_top/la0/la_trig_mask[15] ), 
            .I2(n1865), .O(n1866)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2917.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2918 (.I0(n1866), .I1(n1791), .I2(n1790), .I3(\edb_top/la0/data_out_shift_reg[16] ), 
            .O(n1139)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44 */ ;
    defparam LUT__2918.LUTMASK = 16'h4f44;
    EFX_LUT4 LUT__2919 (.I0(n1779), .I1(\edb_top/la0/la_trig_pos[10] ), 
            .I2(\edb_top/la0/register_conn[66][16] ), .I3(n1777), .O(n1867)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2919.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2920 (.I0(n1792), .I1(\edb_top/la0/register_conn[65][16] ), 
            .I2(n1867), .O(n1868)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2920.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2921 (.I0(n1786), .I1(\edb_top/la0/la_trig_mask[16] ), 
            .I2(n1868), .O(n1869)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2921.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2922 (.I0(n1869), .I1(n1791), .I2(n1790), .I3(\edb_top/la0/data_out_shift_reg[17] ), 
            .O(n1140)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44 */ ;
    defparam LUT__2922.LUTMASK = 16'h4f44;
    EFX_LUT4 LUT__2923 (.I0(n1779), .I1(\edb_top/la0/la_trig_pos[11] ), 
            .I2(\edb_top/la0/register_conn[66][17] ), .I3(n1777), .O(n1870)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2923.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2924 (.I0(n1792), .I1(\edb_top/la0/register_conn[65][17] ), 
            .I2(n1870), .O(n1871)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2924.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2925 (.I0(n1786), .I1(\edb_top/la0/la_trig_mask[17] ), 
            .I2(n1871), .O(n1872)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2925.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2926 (.I0(n1872), .I1(n1791), .I2(n1790), .I3(\edb_top/la0/data_out_shift_reg[18] ), 
            .O(n1141)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44 */ ;
    defparam LUT__2926.LUTMASK = 16'h4f44;
    EFX_LUT4 LUT__2927 (.I0(n1779), .I1(\edb_top/la0/la_trig_pos[12] ), 
            .I2(\edb_top/la0/register_conn[66][18] ), .I3(n1777), .O(n1873)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2927.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2928 (.I0(n1792), .I1(\edb_top/la0/register_conn[65][18] ), 
            .I2(n1873), .O(n1874)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2928.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2929 (.I0(n1786), .I1(\edb_top/la0/la_trig_mask[18] ), 
            .I2(n1874), .O(n1875)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2929.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2930 (.I0(n1875), .I1(n1791), .I2(n1790), .I3(\edb_top/la0/data_out_shift_reg[19] ), 
            .O(n1142)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44 */ ;
    defparam LUT__2930.LUTMASK = 16'h4f44;
    EFX_LUT4 LUT__2931 (.I0(n1779), .I1(\edb_top/la0/la_trig_pos[13] ), 
            .I2(\edb_top/la0/register_conn[66][19] ), .I3(n1777), .O(n1876)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2931.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2932 (.I0(n1792), .I1(\edb_top/la0/register_conn[65][19] ), 
            .I2(n1876), .O(n1877)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2932.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2933 (.I0(n1786), .I1(\edb_top/la0/la_trig_mask[19] ), 
            .I2(n1877), .O(n1878)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2933.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2934 (.I0(n1878), .I1(n1791), .I2(n1790), .I3(\edb_top/la0/data_out_shift_reg[20] ), 
            .O(n1143)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44 */ ;
    defparam LUT__2934.LUTMASK = 16'h4f44;
    EFX_LUT4 LUT__2935 (.I0(n1779), .I1(\edb_top/la0/la_trig_pos[14] ), 
            .I2(\edb_top/la0/register_conn[66][20] ), .I3(n1777), .O(n1879)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2935.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2936 (.I0(n1792), .I1(\edb_top/la0/register_conn[65][20] ), 
            .I2(n1879), .O(n1880)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2936.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2937 (.I0(n1786), .I1(\edb_top/la0/la_trig_mask[20] ), 
            .I2(n1880), .O(n1881)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2937.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2938 (.I0(n1881), .I1(n1791), .I2(n1790), .I3(\edb_top/la0/data_out_shift_reg[21] ), 
            .O(n1144)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44 */ ;
    defparam LUT__2938.LUTMASK = 16'h4f44;
    EFX_LUT4 LUT__2939 (.I0(n1779), .I1(\edb_top/la0/la_trig_pos[15] ), 
            .I2(\edb_top/la0/register_conn[66][21] ), .I3(n1777), .O(n1882)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2939.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2940 (.I0(n1792), .I1(\edb_top/la0/register_conn[65][21] ), 
            .I2(n1882), .O(n1883)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2940.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2941 (.I0(n1786), .I1(\edb_top/la0/la_trig_mask[21] ), 
            .I2(n1883), .O(n1884)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2941.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2942 (.I0(n1884), .I1(n1791), .I2(n1790), .I3(\edb_top/la0/data_out_shift_reg[22] ), 
            .O(n1145)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44 */ ;
    defparam LUT__2942.LUTMASK = 16'h4f44;
    EFX_LUT4 LUT__2943 (.I0(n1779), .I1(\edb_top/la0/la_trig_pos[16] ), 
            .I2(\edb_top/la0/register_conn[66][22] ), .I3(n1777), .O(n1885)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2943.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2944 (.I0(n1792), .I1(\edb_top/la0/register_conn[65][22] ), 
            .I2(n1885), .O(n1886)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2944.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2945 (.I0(n1786), .I1(\edb_top/la0/la_trig_mask[22] ), 
            .I2(n1886), .O(n1887)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2945.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2946 (.I0(n1887), .I1(n1791), .I2(n1790), .I3(\edb_top/la0/data_out_shift_reg[23] ), 
            .O(n1146)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44 */ ;
    defparam LUT__2946.LUTMASK = 16'h4f44;
    EFX_LUT4 LUT__2947 (.I0(n1779), .I1(\edb_top/la0/la_trig_pattern[0] ), 
            .I2(n1777), .I3(\edb_top/la0/register_conn[66][23] ), .O(n1888)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2947.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2948 (.I0(n1792), .I1(\edb_top/la0/register_conn[65][23] ), 
            .I2(n1888), .O(n1889)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2948.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2949 (.I0(n1786), .I1(\edb_top/la0/la_trig_mask[23] ), 
            .I2(n1889), .O(n1890)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2949.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2950 (.I0(n1890), .I1(n1791), .I2(n1790), .I3(\edb_top/la0/data_out_shift_reg[24] ), 
            .O(n1147)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44 */ ;
    defparam LUT__2950.LUTMASK = 16'h4f44;
    EFX_LUT4 LUT__2951 (.I0(n1779), .I1(\edb_top/la0/la_trig_pattern[1] ), 
            .I2(n1777), .I3(\edb_top/la0/register_conn[66][24] ), .O(n1891)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2951.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2952 (.I0(n1792), .I1(\edb_top/la0/register_conn[65][24] ), 
            .I2(n1891), .O(n1892)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2952.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2953 (.I0(n1786), .I1(\edb_top/la0/la_trig_mask[24] ), 
            .I2(n1892), .O(n1893)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2953.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2954 (.I0(n1893), .I1(n1791), .I2(n1790), .I3(\edb_top/la0/data_out_shift_reg[25] ), 
            .O(n1148)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44 */ ;
    defparam LUT__2954.LUTMASK = 16'h4f44;
    EFX_LUT4 LUT__2955 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][25] ), 
            .I2(\edb_top/la0/la_trig_mask[25] ), .I3(n1786), .O(n1894)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2955.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2956 (.I0(\edb_top/la0/register_conn[65][25] ), .I1(n1792), 
            .I2(n1894), .I3(n1791), .O(n1895)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__2956.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__2957 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[26] ), 
            .I2(n1895), .O(n1149)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__2957.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__2958 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][26] ), 
            .I2(\edb_top/la0/la_trig_mask[26] ), .I3(n1786), .O(n1896)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2958.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2959 (.I0(\edb_top/la0/register_conn[65][26] ), .I1(n1792), 
            .I2(n1896), .I3(n1791), .O(n1897)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__2959.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__2960 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[27] ), 
            .I2(n1897), .O(n1150)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__2960.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__2961 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][27] ), 
            .I2(\edb_top/la0/la_trig_mask[27] ), .I3(n1786), .O(n1898)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2961.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2962 (.I0(\edb_top/la0/register_conn[65][27] ), .I1(n1792), 
            .I2(n1898), .I3(n1791), .O(n1899)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__2962.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__2963 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[28] ), 
            .I2(n1899), .O(n1151)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__2963.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__2964 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][28] ), 
            .I2(\edb_top/la0/la_trig_mask[28] ), .I3(n1786), .O(n1900)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2964.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2965 (.I0(\edb_top/la0/register_conn[65][28] ), .I1(n1792), 
            .I2(n1900), .I3(n1791), .O(n1901)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__2965.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__2966 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[29] ), 
            .I2(n1901), .O(n1152)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__2966.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__2967 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][29] ), 
            .I2(\edb_top/la0/la_trig_mask[29] ), .I3(n1786), .O(n1902)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2967.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2968 (.I0(\edb_top/la0/register_conn[65][29] ), .I1(n1792), 
            .I2(n1902), .I3(n1791), .O(n1903)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__2968.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__2969 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[30] ), 
            .I2(n1903), .O(n1153)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__2969.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__2970 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][30] ), 
            .I2(\edb_top/la0/la_trig_mask[30] ), .I3(n1786), .O(n1904)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2970.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2971 (.I0(\edb_top/la0/register_conn[65][30] ), .I1(n1792), 
            .I2(n1904), .I3(n1791), .O(n1905)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__2971.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__2972 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[31] ), 
            .I2(n1905), .O(n1154)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__2972.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__2973 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][31] ), 
            .I2(\edb_top/la0/la_trig_mask[31] ), .I3(n1786), .O(n1906)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2973.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2974 (.I0(\edb_top/la0/register_conn[65][31] ), .I1(n1792), 
            .I2(n1906), .I3(n1791), .O(n1907)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__2974.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__2975 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[32] ), 
            .I2(n1907), .O(n1155)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__2975.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__2976 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][32] ), 
            .I2(\edb_top/la0/la_trig_mask[32] ), .I3(n1786), .O(n1908)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2976.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2977 (.I0(\edb_top/la0/register_conn[65][32] ), .I1(n1792), 
            .I2(n1908), .I3(n1791), .O(n1909)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__2977.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__2978 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[33] ), 
            .I2(n1909), .O(n1156)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__2978.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__2979 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][33] ), 
            .I2(\edb_top/la0/la_trig_mask[33] ), .I3(n1786), .O(n1910)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2979.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2980 (.I0(\edb_top/la0/register_conn[65][33] ), .I1(n1792), 
            .I2(n1910), .I3(n1791), .O(n1911)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__2980.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__2981 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[34] ), 
            .I2(n1911), .O(n1157)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__2981.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__2982 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][34] ), 
            .I2(\edb_top/la0/la_trig_mask[34] ), .I3(n1786), .O(n1912)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2982.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2983 (.I0(\edb_top/la0/register_conn[65][34] ), .I1(n1792), 
            .I2(n1912), .I3(n1791), .O(n1913)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__2983.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__2984 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[35] ), 
            .I2(n1913), .O(n1158)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__2984.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__2985 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][35] ), 
            .I2(\edb_top/la0/la_trig_mask[35] ), .I3(n1786), .O(n1914)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2985.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2986 (.I0(\edb_top/la0/register_conn[65][35] ), .I1(n1792), 
            .I2(n1914), .I3(n1791), .O(n1915)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__2986.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__2987 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[36] ), 
            .I2(n1915), .O(n1159)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__2987.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__2988 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][36] ), 
            .I2(\edb_top/la0/la_trig_mask[36] ), .I3(n1786), .O(n1916)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2988.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2989 (.I0(\edb_top/la0/register_conn[65][36] ), .I1(n1792), 
            .I2(n1916), .I3(n1791), .O(n1917)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__2989.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__2990 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[37] ), 
            .I2(n1917), .O(n1160)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__2990.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__2991 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][37] ), 
            .I2(\edb_top/la0/la_trig_mask[37] ), .I3(n1786), .O(n1918)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2991.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2992 (.I0(\edb_top/la0/register_conn[65][37] ), .I1(n1792), 
            .I2(n1918), .I3(n1791), .O(n1919)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__2992.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__2993 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[38] ), 
            .I2(n1919), .O(n1161)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__2993.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__2994 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][38] ), 
            .I2(\edb_top/la0/la_trig_mask[38] ), .I3(n1786), .O(n1920)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2994.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2995 (.I0(\edb_top/la0/register_conn[65][38] ), .I1(n1792), 
            .I2(n1920), .I3(n1791), .O(n1921)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__2995.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__2996 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[39] ), 
            .I2(n1921), .O(n1162)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__2996.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__2997 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][39] ), 
            .I2(\edb_top/la0/la_trig_mask[39] ), .I3(n1786), .O(n1922)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2997.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2998 (.I0(\edb_top/la0/register_conn[65][39] ), .I1(n1792), 
            .I2(n1922), .I3(n1791), .O(n1923)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__2998.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__2999 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[40] ), 
            .I2(n1923), .O(n1163)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__2999.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__3000 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][40] ), 
            .I2(\edb_top/la0/la_trig_mask[40] ), .I3(n1786), .O(n1924)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3000.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3001 (.I0(\edb_top/la0/register_conn[65][40] ), .I1(n1792), 
            .I2(n1924), .I3(n1791), .O(n1925)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__3001.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__3002 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[41] ), 
            .I2(n1925), .O(n1164)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__3002.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__3003 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][41] ), 
            .I2(\edb_top/la0/la_trig_mask[41] ), .I3(n1786), .O(n1926)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3003.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3004 (.I0(\edb_top/la0/register_conn[65][41] ), .I1(n1792), 
            .I2(n1926), .I3(n1791), .O(n1927)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__3004.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__3005 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[42] ), 
            .I2(n1927), .O(n1165)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__3005.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__3006 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][42] ), 
            .I2(\edb_top/la0/la_trig_mask[42] ), .I3(n1786), .O(n1928)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3006.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3007 (.I0(\edb_top/la0/register_conn[65][42] ), .I1(n1792), 
            .I2(n1928), .I3(n1791), .O(n1929)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__3007.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__3008 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[43] ), 
            .I2(n1929), .O(n1166)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__3008.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__3009 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][43] ), 
            .I2(\edb_top/la0/la_trig_mask[43] ), .I3(n1786), .O(n1930)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3009.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3010 (.I0(\edb_top/la0/register_conn[65][43] ), .I1(n1792), 
            .I2(n1930), .I3(n1791), .O(n1931)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__3010.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__3011 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[44] ), 
            .I2(n1931), .O(n1167)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__3011.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__3012 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][44] ), 
            .I2(\edb_top/la0/la_trig_mask[44] ), .I3(n1786), .O(n1932)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3012.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3013 (.I0(\edb_top/la0/register_conn[65][44] ), .I1(n1792), 
            .I2(n1932), .I3(n1791), .O(n1933)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__3013.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__3014 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[45] ), 
            .I2(n1933), .O(n1168)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__3014.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__3015 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][45] ), 
            .I2(\edb_top/la0/la_trig_mask[45] ), .I3(n1786), .O(n1934)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3015.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3016 (.I0(\edb_top/la0/register_conn[65][45] ), .I1(n1792), 
            .I2(n1934), .I3(n1791), .O(n1935)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__3016.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__3017 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[46] ), 
            .I2(n1935), .O(n1169)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__3017.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__3018 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][46] ), 
            .I2(\edb_top/la0/la_trig_mask[46] ), .I3(n1786), .O(n1936)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3018.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3019 (.I0(\edb_top/la0/register_conn[65][46] ), .I1(n1792), 
            .I2(n1936), .I3(n1791), .O(n1937)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__3019.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__3020 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[47] ), 
            .I2(n1937), .O(n1170)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__3020.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__3021 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][47] ), 
            .I2(\edb_top/la0/la_trig_mask[47] ), .I3(n1786), .O(n1938)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3021.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3022 (.I0(\edb_top/la0/register_conn[65][47] ), .I1(n1792), 
            .I2(n1938), .I3(n1791), .O(n1939)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__3022.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__3023 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[48] ), 
            .I2(n1939), .O(n1171)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__3023.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__3024 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][48] ), 
            .I2(\edb_top/la0/la_trig_mask[48] ), .I3(n1786), .O(n1940)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3024.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3025 (.I0(\edb_top/la0/register_conn[65][48] ), .I1(n1792), 
            .I2(n1940), .I3(n1791), .O(n1941)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__3025.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__3026 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[49] ), 
            .I2(n1941), .O(n1172)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__3026.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__3027 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][49] ), 
            .I2(\edb_top/la0/la_trig_mask[49] ), .I3(n1786), .O(n1942)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3027.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3028 (.I0(\edb_top/la0/register_conn[65][49] ), .I1(n1792), 
            .I2(n1942), .I3(n1791), .O(n1943)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__3028.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__3029 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[50] ), 
            .I2(n1943), .O(n1173)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__3029.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__3030 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][50] ), 
            .I2(\edb_top/la0/la_trig_mask[50] ), .I3(n1786), .O(n1944)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3030.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3031 (.I0(\edb_top/la0/register_conn[65][50] ), .I1(n1792), 
            .I2(n1944), .I3(n1791), .O(n1945)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__3031.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__3032 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[51] ), 
            .I2(n1945), .O(n1174)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__3032.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__3033 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][51] ), 
            .I2(\edb_top/la0/la_trig_mask[51] ), .I3(n1786), .O(n1946)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3033.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3034 (.I0(\edb_top/la0/register_conn[65][51] ), .I1(n1792), 
            .I2(n1946), .I3(n1791), .O(n1947)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__3034.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__3035 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[52] ), 
            .I2(n1947), .O(n1175)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__3035.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__3036 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][52] ), 
            .I2(\edb_top/la0/la_trig_mask[52] ), .I3(n1786), .O(n1948)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3036.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3037 (.I0(\edb_top/la0/register_conn[65][52] ), .I1(n1792), 
            .I2(n1948), .I3(n1791), .O(n1949)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__3037.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__3038 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[53] ), 
            .I2(n1949), .O(n1176)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__3038.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__3039 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][53] ), 
            .I2(\edb_top/la0/la_trig_mask[53] ), .I3(n1786), .O(n1950)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3039.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3040 (.I0(\edb_top/la0/register_conn[65][53] ), .I1(n1792), 
            .I2(n1950), .I3(n1791), .O(n1951)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__3040.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__3041 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[54] ), 
            .I2(n1951), .O(n1177)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__3041.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__3042 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][54] ), 
            .I2(\edb_top/la0/la_trig_mask[54] ), .I3(n1786), .O(n1952)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3042.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3043 (.I0(\edb_top/la0/register_conn[65][54] ), .I1(n1792), 
            .I2(n1952), .I3(n1791), .O(n1953)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__3043.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__3044 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[55] ), 
            .I2(n1953), .O(n1178)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__3044.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__3045 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][55] ), 
            .I2(\edb_top/la0/la_trig_mask[55] ), .I3(n1786), .O(n1954)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3045.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3046 (.I0(\edb_top/la0/register_conn[65][55] ), .I1(n1792), 
            .I2(n1954), .I3(n1791), .O(n1955)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__3046.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__3047 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[56] ), 
            .I2(n1955), .O(n1179)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__3047.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__3048 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][56] ), 
            .I2(\edb_top/la0/la_trig_mask[56] ), .I3(n1786), .O(n1956)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3048.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3049 (.I0(\edb_top/la0/register_conn[65][56] ), .I1(n1792), 
            .I2(n1956), .I3(n1791), .O(n1957)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__3049.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__3050 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[57] ), 
            .I2(n1957), .O(n1180)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__3050.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__3051 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][57] ), 
            .I2(\edb_top/la0/la_trig_mask[57] ), .I3(n1786), .O(n1958)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3051.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3052 (.I0(\edb_top/la0/register_conn[65][57] ), .I1(n1792), 
            .I2(n1958), .I3(n1791), .O(n1959)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__3052.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__3053 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[58] ), 
            .I2(n1959), .O(n1181)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__3053.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__3054 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][58] ), 
            .I2(\edb_top/la0/la_trig_mask[58] ), .I3(n1786), .O(n1960)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3054.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3055 (.I0(\edb_top/la0/register_conn[65][58] ), .I1(n1792), 
            .I2(n1960), .I3(n1791), .O(n1961)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__3055.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__3056 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[59] ), 
            .I2(n1961), .O(n1182)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__3056.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__3057 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][59] ), 
            .I2(\edb_top/la0/la_trig_mask[59] ), .I3(n1786), .O(n1962)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3057.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3058 (.I0(\edb_top/la0/register_conn[65][59] ), .I1(n1792), 
            .I2(n1962), .I3(n1791), .O(n1963)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__3058.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__3059 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[60] ), 
            .I2(n1963), .O(n1183)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__3059.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__3060 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][60] ), 
            .I2(\edb_top/la0/la_trig_mask[60] ), .I3(n1786), .O(n1964)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3060.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3061 (.I0(\edb_top/la0/register_conn[65][60] ), .I1(n1792), 
            .I2(n1964), .I3(n1791), .O(n1965)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__3061.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__3062 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[61] ), 
            .I2(n1965), .O(n1184)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__3062.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__3063 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][61] ), 
            .I2(\edb_top/la0/la_trig_mask[61] ), .I3(n1786), .O(n1966)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3063.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3064 (.I0(\edb_top/la0/register_conn[65][61] ), .I1(n1792), 
            .I2(n1966), .I3(n1791), .O(n1967)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__3064.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__3065 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[62] ), 
            .I2(n1967), .O(n1185)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__3065.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__3066 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][62] ), 
            .I2(\edb_top/la0/la_trig_mask[62] ), .I3(n1786), .O(n1968)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3066.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3067 (.I0(\edb_top/la0/register_conn[65][62] ), .I1(n1792), 
            .I2(n1968), .I3(n1791), .O(n1969)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__3067.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__3068 (.I0(n1790), .I1(\edb_top/la0/data_out_shift_reg[63] ), 
            .I2(n1969), .O(n1186)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__3068.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__3069 (.I0(n1777), .I1(\edb_top/la0/register_conn[66][63] ), 
            .I2(\edb_top/la0/la_trig_mask[63] ), .I3(n1786), .O(n1970)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3069.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3070 (.I0(\edb_top/la0/register_conn[65][63] ), .I1(n1792), 
            .I2(n1970), .I3(n1791), .O(n1187)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__3070.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__3071 (.I0(n1684), .I1(\edb_top/la0/module_state[2] ), 
            .I2(\edb_top/la0/module_state[3] ), .I3(n1738), .O(n1971)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__3071.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__3072 (.I0(bscan_UPDATE), .I1(n1753), .I2(\edb_top/la0/module_state[1] ), 
            .O(n1972)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3072.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3073 (.I0(bscan_UPDATE), .I1(\edb_top/la0/module_state[1] ), 
            .I2(\edb_top/la0/module_state[0] ), .I3(\edb_top/la0/module_state[3] ), 
            .O(n1973)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h050c */ ;
    defparam LUT__3073.LUTMASK = 16'h050c;
    EFX_LUT4 LUT__3074 (.I0(n1686), .I1(n1973), .I2(\edb_top/la0/module_state[2] ), 
            .I3(n1972), .O(n1974)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f1 */ ;
    defparam LUT__3074.LUTMASK = 16'h00f1;
    EFX_LUT4 LUT__3075 (.I0(n1697), .I1(n1971), .I2(n1974), .O(n1188)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f4f */ ;
    defparam LUT__3075.LUTMASK = 16'h4f4f;
    EFX_LUT4 LUT__3076 (.I0(n1761), .I1(n1764), .I2(n1765), .O(n1975)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__3076.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__3077 (.I0(n1752), .I1(\edb_top/la0/module_state[0] ), 
            .I2(\edb_top/la0/module_state[1] ), .O(n1976)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171 */ ;
    defparam LUT__3077.LUTMASK = 16'h7171;
    EFX_LUT4 LUT__3078 (.I0(bscan_UPDATE), .I1(n1976), .I2(n1753), .I3(n1762), 
            .O(n1977)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf */ ;
    defparam LUT__3078.LUTMASK = 16'h00bf;
    EFX_LUT4 LUT__3079 (.I0(n1738), .I1(bscan_UPDATE), .I2(n1697), .O(n1978)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__3079.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__3080 (.I0(n1753), .I1(n1975), .I2(n1978), .I3(n1977), 
            .O(n1189)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0ff */ ;
    defparam LUT__3080.LUTMASK = 16'he0ff;
    EFX_LUT4 LUT__3081 (.I0(n1754), .I1(n1765), .I2(n1699), .I3(n1697), 
            .O(n1979)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfa30 */ ;
    defparam LUT__3081.LUTMASK = 16'hfa30;
    EFX_LUT4 LUT__3082 (.I0(bscan_UPDATE), .I1(n1979), .O(n1190)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3082.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3083 (.I0(n990), .I1(\edb_top/la0/crc_data_out[1] ), .O(n1191)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__3083.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__3084 (.I0(n990), .I1(n1771), .I2(n1277), .O(n1192)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__3084.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__3085 (.I0(n990), .I1(\edb_top/la0/crc_data_out[2] ), .O(n1193)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__3085.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__3086 (.I0(n990), .I1(\edb_top/la0/crc_data_out[3] ), .O(n1194)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__3086.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__3087 (.I0(n990), .I1(\edb_top/la0/crc_data_out[4] ), .O(n1195)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__3087.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__3088 (.I0(n990), .I1(\edb_top/la0/crc_data_out[5] ), .O(n1196)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__3088.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__3089 (.I0(bscan_TDI), .I1(\edb_top/la0/data_out_shift_reg[0] ), 
            .I2(\edb_top/la0/module_state[1] ), .I3(\edb_top/la0/crc_data_out[0] ), 
            .O(n1980)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac53 */ ;
    defparam LUT__3089.LUTMASK = 16'hac53;
    EFX_LUT4 LUT__3090 (.I0(n1980), .I1(n1771), .O(n1981)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3090.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3091 (.I0(n990), .I1(n1981), .I2(\edb_top/la0/crc_data_out[6] ), 
            .O(n1197)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e */ ;
    defparam LUT__3091.LUTMASK = 16'h3e3e;
    EFX_LUT4 LUT__3092 (.I0(n990), .I1(\edb_top/la0/crc_data_out[7] ), .O(n1199)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__3092.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__3093 (.I0(n990), .I1(\edb_top/la0/crc_data_out[8] ), .O(n1200)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__3093.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__3094 (.I0(n990), .I1(n1981), .I2(\edb_top/la0/crc_data_out[9] ), 
            .O(n1201)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e */ ;
    defparam LUT__3094.LUTMASK = 16'h3e3e;
    EFX_LUT4 LUT__3095 (.I0(n990), .I1(n1981), .I2(\edb_top/la0/crc_data_out[10] ), 
            .O(n1202)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e */ ;
    defparam LUT__3095.LUTMASK = 16'h3e3e;
    EFX_LUT4 LUT__3096 (.I0(n990), .I1(\edb_top/la0/crc_data_out[11] ), 
            .O(n1203)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__3096.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__3097 (.I0(n990), .I1(\edb_top/la0/crc_data_out[12] ), 
            .O(n1204)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__3097.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__3098 (.I0(n990), .I1(\edb_top/la0/crc_data_out[13] ), 
            .O(n1205)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__3098.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__3099 (.I0(n990), .I1(\edb_top/la0/crc_data_out[14] ), 
            .O(n1206)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__3099.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__3100 (.I0(n990), .I1(\edb_top/la0/crc_data_out[15] ), 
            .O(n1207)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__3100.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__3101 (.I0(n990), .I1(n1981), .I2(\edb_top/la0/crc_data_out[16] ), 
            .O(n1208)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e */ ;
    defparam LUT__3101.LUTMASK = 16'h3e3e;
    EFX_LUT4 LUT__3102 (.I0(n990), .I1(\edb_top/la0/crc_data_out[17] ), 
            .O(n1209)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__3102.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__3103 (.I0(n990), .I1(\edb_top/la0/crc_data_out[18] ), 
            .O(n1210)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__3103.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__3104 (.I0(n990), .I1(\edb_top/la0/crc_data_out[19] ), 
            .O(n1211)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__3104.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__3105 (.I0(n990), .I1(n1981), .I2(\edb_top/la0/crc_data_out[20] ), 
            .O(n1212)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e */ ;
    defparam LUT__3105.LUTMASK = 16'h3e3e;
    EFX_LUT4 LUT__3106 (.I0(n990), .I1(n1981), .I2(\edb_top/la0/crc_data_out[21] ), 
            .O(n1213)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e */ ;
    defparam LUT__3106.LUTMASK = 16'h3e3e;
    EFX_LUT4 LUT__3107 (.I0(n990), .I1(n1981), .I2(\edb_top/la0/crc_data_out[22] ), 
            .O(n1214)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e */ ;
    defparam LUT__3107.LUTMASK = 16'h3e3e;
    EFX_LUT4 LUT__3108 (.I0(n990), .I1(\edb_top/la0/crc_data_out[23] ), 
            .O(n1215)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__3108.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__3109 (.I0(n990), .I1(n1981), .I2(\edb_top/la0/crc_data_out[24] ), 
            .O(n1216)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e */ ;
    defparam LUT__3109.LUTMASK = 16'h3e3e;
    EFX_LUT4 LUT__3110 (.I0(n990), .I1(n1981), .I2(\edb_top/la0/crc_data_out[25] ), 
            .O(n1217)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e */ ;
    defparam LUT__3110.LUTMASK = 16'h3e3e;
    EFX_LUT4 LUT__3111 (.I0(n990), .I1(\edb_top/la0/crc_data_out[26] ), 
            .O(n1218)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__3111.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__3112 (.I0(n990), .I1(n1981), .I2(\edb_top/la0/crc_data_out[27] ), 
            .O(n1219)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e */ ;
    defparam LUT__3112.LUTMASK = 16'h3e3e;
    EFX_LUT4 LUT__3113 (.I0(n990), .I1(n1981), .I2(\edb_top/la0/crc_data_out[28] ), 
            .O(n1220)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e */ ;
    defparam LUT__3113.LUTMASK = 16'h3e3e;
    EFX_LUT4 LUT__3114 (.I0(n990), .I1(\edb_top/la0/crc_data_out[29] ), 
            .O(n1221)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__3114.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__3115 (.I0(n990), .I1(n1981), .I2(\edb_top/la0/crc_data_out[30] ), 
            .O(n1222)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e */ ;
    defparam LUT__3115.LUTMASK = 16'h3e3e;
    EFX_LUT4 LUT__3116 (.I0(n990), .I1(n1981), .I2(\edb_top/la0/crc_data_out[31] ), 
            .O(n1223)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e */ ;
    defparam LUT__3116.LUTMASK = 16'h3e3e;
    EFX_LUT4 LUT__3117 (.I0(n1981), .I1(n990), .O(n1224)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__3117.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__3118 (.I0(\edb_top/la0/register_conn[65][0] ), .I1(\edb_top/la0/register_conn[66][0] ), 
            .O(n1239)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3118.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3119 (.I0(\edb_top/la0/cap_fifo_din[5] ), .I1(\edb_top/la0/register_conn[65][5] ), 
            .I2(\edb_top/la0/cap_fifo_din[6] ), .I3(\edb_top/la0/register_conn[65][6] ), 
            .O(n1982)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__3119.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__3120 (.I0(\edb_top/la0/cap_fifo_din[4] ), .I1(\edb_top/la0/register_conn[65][4] ), 
            .I2(\edb_top/la0/cap_fifo_din[7] ), .I3(\edb_top/la0/register_conn[65][7] ), 
            .O(n1983)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__3120.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__3121 (.I0(n1982), .I1(n1983), .O(n1984)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3121.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3122 (.I0(\edb_top/la0/cap_fifo_din[3] ), .I1(\edb_top/la0/register_conn[65][3] ), 
            .I2(\edb_top/la0/register_conn[65][2] ), .I3(\edb_top/la0/cap_fifo_din[2] ), 
            .O(n1985)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__3122.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__3123 (.I0(\edb_top/la0/register_conn[65][4] ), .I1(\edb_top/la0/cap_fifo_din[4] ), 
            .I2(n1985), .I3(n1984), .O(n1986)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__3123.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__3124 (.I0(\edb_top/la0/cap_fifo_din[6] ), .I1(\edb_top/la0/register_conn[65][6] ), 
            .I2(\edb_top/la0/register_conn[65][5] ), .I3(\edb_top/la0/cap_fifo_din[5] ), 
            .O(n1987)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__3124.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__3125 (.I0(n1987), .I1(\edb_top/la0/cap_fifo_din[7] ), 
            .I2(\edb_top/la0/register_conn[65][7] ), .I3(n1986), .O(n1988)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2 */ ;
    defparam LUT__3125.LUTMASK = 16'h00b2;
    EFX_LUT4 LUT__3126 (.I0(\edb_top/la0/cap_fifo_din[1] ), .I1(\edb_top/la0/register_conn[65][1] ), 
            .I2(\edb_top/la0/cap_fifo_din[2] ), .I3(\edb_top/la0/register_conn[65][2] ), 
            .O(n1989)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__3126.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__3127 (.I0(\edb_top/la0/cap_fifo_din[3] ), .I1(\edb_top/la0/register_conn[65][3] ), 
            .I2(n1984), .I3(n1989), .O(n1990)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb000 */ ;
    defparam LUT__3127.LUTMASK = 16'hb000;
    EFX_LUT4 LUT__3128 (.I0(\edb_top/la0/cap_fifo_din[1] ), .I1(\edb_top/la0/register_conn[65][1] ), 
            .I2(\edb_top/la0/cap_fifo_din[0] ), .I3(\edb_top/la0/register_conn[65][0] ), 
            .O(n1991)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__3128.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__3129 (.I0(n1990), .I1(n1991), .I2(n1988), .O(n1240)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__3129.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__3130 (.I0(\edb_top/la0/register_conn[65][0] ), .I1(\edb_top/la0/cap_fifo_din[0] ), 
            .I2(\edb_top/la0/register_conn[65][1] ), .I3(\edb_top/la0/cap_fifo_din[1] ), 
            .O(n1992)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__3130.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__3131 (.I0(n1990), .I1(n1992), .I2(n1988), .O(n1241)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__3131.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__3132 (.I0(\edb_top/la0/cap_fifo_din[0] ), .I1(\edb_top/la0/register_conn[66][0] ), 
            .O(n1242)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3132.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3133 (.I0(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[4] ), 
            .I1(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[4] ), .I2(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[7] ), 
            .I3(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[7] ), .O(n1993)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__3133.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__3134 (.I0(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[2] ), 
            .I1(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[2] ), .I2(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[3] ), 
            .I3(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[3] ), .O(n1994)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__3134.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__3135 (.I0(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[0] ), 
            .I1(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[0] ), .I2(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[1] ), 
            .I3(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[1] ), .O(n1995)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__3135.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__3136 (.I0(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[5] ), 
            .I1(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[5] ), .I2(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp2[6] ), 
            .I3(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp1[6] ), .O(n1996)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__3136.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__3137 (.I0(n1993), .I1(n1994), .I2(n1995), .I3(n1996), 
            .O(n1997)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__3137.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__3138 (.I0(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp3[0] ), 
            .I1(n1997), .I2(\edb_top/la0/register_conn[64][0] ), .I3(\edb_top/la0/register_conn[64][1] ), 
            .O(n1998)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3c0 */ ;
    defparam LUT__3138.LUTMASK = 16'ha3c0;
    EFX_LUT4 LUT__3139 (.I0(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp6[0] ), 
            .I1(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp4[0] ), .I2(\edb_top/la0/register_conn[64][1] ), 
            .O(n1999)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__3139.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__3140 (.I0(\edb_top/la0/register_conn[64][1] ), .I1(\edb_top/la0/GEN_PROBE[0].compare_unit_inst/exp5[0] ), 
            .I2(n1999), .I3(\edb_top/la0/register_conn[64][0] ), .O(n2000)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__3140.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__3141 (.I0(n1998), .I1(n2000), .I2(\edb_top/la0/register_conn[64][2] ), 
            .O(n1243)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__3141.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__3142 (.I0(\edb_top/la0/register_conn[65][1] ), .I1(\edb_top/la0/register_conn[66][1] ), 
            .O(n1244)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3142.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3143 (.I0(\edb_top/la0/register_conn[65][2] ), .I1(\edb_top/la0/register_conn[66][2] ), 
            .O(n1245)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3143.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3144 (.I0(\edb_top/la0/register_conn[65][3] ), .I1(\edb_top/la0/register_conn[66][3] ), 
            .O(n1246)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3144.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3145 (.I0(\edb_top/la0/register_conn[65][4] ), .I1(\edb_top/la0/register_conn[66][4] ), 
            .O(n1247)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3145.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3146 (.I0(\edb_top/la0/register_conn[65][5] ), .I1(\edb_top/la0/register_conn[66][5] ), 
            .O(n1248)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3146.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3147 (.I0(\edb_top/la0/register_conn[65][6] ), .I1(\edb_top/la0/register_conn[66][6] ), 
            .O(n1249)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3147.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3148 (.I0(\edb_top/la0/register_conn[65][7] ), .I1(\edb_top/la0/register_conn[66][7] ), 
            .O(n1250)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3148.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3149 (.I0(\edb_top/la0/cap_fifo_din[1] ), .I1(\edb_top/la0/register_conn[66][1] ), 
            .O(n1251)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3149.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3150 (.I0(\edb_top/la0/cap_fifo_din[2] ), .I1(\edb_top/la0/register_conn[66][2] ), 
            .O(n1252)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3150.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3151 (.I0(\edb_top/la0/cap_fifo_din[3] ), .I1(\edb_top/la0/register_conn[66][3] ), 
            .O(n1253)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3151.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3152 (.I0(\edb_top/la0/cap_fifo_din[4] ), .I1(\edb_top/la0/register_conn[66][4] ), 
            .O(n1254)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3152.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3153 (.I0(\edb_top/la0/cap_fifo_din[5] ), .I1(\edb_top/la0/register_conn[66][5] ), 
            .O(n1255)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3153.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3154 (.I0(\edb_top/la0/cap_fifo_din[6] ), .I1(\edb_top/la0/register_conn[66][6] ), 
            .O(n1256)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3154.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3155 (.I0(\edb_top/la0/cap_fifo_din[7] ), .I1(\edb_top/la0/register_conn[66][7] ), 
            .O(n1257)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3155.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3156 (.I0(\edb_top/la0/la_trig_pattern[1] ), .I1(\edb_top/la0/tu_data[0] ), 
            .I2(\edb_top/la0/la_trig_mask[0] ), .O(n1258)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__3156.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__3157 (.I0(\edb_top/la0/la_biu_inst/cap_buf_read_done_p2 ), 
            .I1(n635), .O(n1282)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3157.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3158 (.I0(\edb_top/la0/register_conn[0][2] ), .I1(\edb_top/la0/register_conn[0][1] ), 
            .I2(\edb_top/la0/register_conn[0][0] ), .I3(\edb_top/la0/la_biu_inst/cap_buf_read_done_p2 ), 
            .O(n1283)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__3158.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__3159 (.I0(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2] ), 
            .I1(\edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]_2 ), 
            .I2(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3] ), 
            .I3(\edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]_2 ), 
            .O(n2001)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__3159.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__3160 (.I0(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6] ), 
            .I1(\edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]_2 ), 
            .I2(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7] ), 
            .I3(\edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]_2 ), 
            .O(n2002)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__3160.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__3161 (.I0(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4] ), 
            .I1(\edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]_2 ), 
            .I2(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5] ), 
            .I3(\edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]_2 ), 
            .O(n2003)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__3161.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__3162 (.I0(n2001), .I1(n2002), .I2(n2003), .O(n2004)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__3162.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__3163 (.I0(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8] ), 
            .I1(\edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]_2 ), 
            .I2(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9] ), 
            .I3(\edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]_2 ), 
            .O(n2005)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__3163.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__3164 (.I0(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0] ), 
            .I1(\edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]_2 ), 
            .I2(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1] ), 
            .I3(\edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]_2 ), 
            .O(n2006)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__3164.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__3165 (.I0(n2004), .I1(n2005), .I2(n2006), .O(n2007)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__3165.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__3166 (.I0(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10] ), 
            .I1(\edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] ), 
            .I2(n2007), .O(n2008)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__3166.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__3167 (.I0(\edb_top/la0/register_conn[0][0] ), .I1(\edb_top/la0/tu_trigger ), 
            .I2(\edb_top/la0/la_biu_inst/run_trig_imdt_p2 ), .I3(\edb_top/la0/register_conn[0][1] ), 
            .O(n2009)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__3167.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__3168 (.I0(n2008), .I1(\edb_top/la0/register_conn[0][0] ), 
            .I2(n2009), .O(n2010)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__3168.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__3169 (.I0(\edb_top/la0/la_biu_inst/pos_counter[9] ), .I1(\edb_top/la0/la_trig_pos[9] ), 
            .I2(\edb_top/la0/register_conn[0][0] ), .O(n2011)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090 */ ;
    defparam LUT__3169.LUTMASK = 16'h9090;
    EFX_LUT4 LUT__3170 (.I0(\edb_top/la0/la_biu_inst/pos_counter[2] ), .I1(\edb_top/la0/la_trig_pos[2] ), 
            .I2(\edb_top/la0/la_biu_inst/pos_counter[11] ), .I3(\edb_top/la0/la_trig_pos[11] ), 
            .O(n2012)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__3170.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__3171 (.I0(\edb_top/la0/la_biu_inst/pos_counter[6] ), .I1(\edb_top/la0/la_trig_pos[6] ), 
            .I2(\edb_top/la0/la_trig_pos[5] ), .I3(\edb_top/la0/la_biu_inst/pos_counter[5] ), 
            .O(n2013)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__3171.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__3172 (.I0(n2011), .I1(n2012), .I2(n2013), .O(n2014)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__3172.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__3173 (.I0(\edb_top/la0/la_biu_inst/pos_counter[13] ), .I1(\edb_top/la0/la_trig_pos[13] ), 
            .I2(\edb_top/la0/la_trig_pos[3] ), .I3(\edb_top/la0/la_biu_inst/pos_counter[3] ), 
            .O(n2015)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__3173.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__3174 (.I0(\edb_top/la0/la_biu_inst/pos_counter[1] ), .I1(\edb_top/la0/la_trig_pos[1] ), 
            .I2(\edb_top/la0/la_biu_inst/pos_counter[16] ), .I3(\edb_top/la0/la_trig_pos[16] ), 
            .O(n2016)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__3174.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__3175 (.I0(\edb_top/la0/la_biu_inst/pos_counter[15] ), .I1(\edb_top/la0/la_trig_pos[15] ), 
            .I2(\edb_top/la0/la_trig_pos[4] ), .I3(\edb_top/la0/la_biu_inst/pos_counter[4] ), 
            .O(n2017)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__3175.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__3176 (.I0(\edb_top/la0/la_biu_inst/pos_counter[10] ), .I1(\edb_top/la0/la_trig_pos[10] ), 
            .I2(\edb_top/la0/la_trig_pos[7] ), .I3(\edb_top/la0/la_biu_inst/pos_counter[7] ), 
            .O(n2018)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__3176.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__3177 (.I0(n2015), .I1(n2016), .I2(n2017), .I3(n2018), 
            .O(n2019)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__3177.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__3178 (.I0(\edb_top/la0/la_biu_inst/pos_counter[12] ), .I1(\edb_top/la0/la_trig_pos[12] ), 
            .I2(\edb_top/la0/la_trig_pos[8] ), .I3(\edb_top/la0/la_biu_inst/pos_counter[8] ), 
            .O(n2020)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__3178.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__3179 (.I0(\edb_top/la0/la_trig_pos[0] ), .I1(\edb_top/la0/la_biu_inst/pos_counter[0] ), 
            .I2(\edb_top/la0/la_biu_inst/pos_counter[14] ), .I3(\edb_top/la0/la_trig_pos[14] ), 
            .O(n2021)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__3179.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__3180 (.I0(n2014), .I1(n2019), .I2(n2020), .I3(n2021), 
            .O(n2022)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__3180.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__3181 (.I0(n2022), .I1(\edb_top/la0/register_conn[0][1] ), 
            .O(n2023)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__3181.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__3182 (.I0(\edb_top/la0/la_trig_pos[13] ), .I1(\edb_top/la0/la_trig_pos[14] ), 
            .I2(\edb_top/la0/la_trig_pos[15] ), .O(n2024)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__3182.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__3183 (.I0(\edb_top/la0/la_trig_pos[9] ), .I1(\edb_top/la0/la_trig_pos[10] ), 
            .I2(\edb_top/la0/la_trig_pos[11] ), .I3(\edb_top/la0/la_trig_pos[12] ), 
            .O(n2025)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3183.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3184 (.I0(\edb_top/la0/la_trig_pos[5] ), .I1(\edb_top/la0/la_trig_pos[6] ), 
            .I2(\edb_top/la0/la_trig_pos[8] ), .I3(\edb_top/la0/la_trig_pos[16] ), 
            .O(n2026)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3184.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3185 (.I0(n2024), .I1(n2025), .I2(n2026), .O(n2027)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__3185.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__3186 (.I0(\edb_top/la0/la_trig_pos[1] ), .I1(\edb_top/la0/la_trig_pos[2] ), 
            .I2(\edb_top/la0/la_trig_pos[3] ), .I3(\edb_top/la0/la_trig_pos[4] ), 
            .O(n2028)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3186.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3187 (.I0(\edb_top/la0/la_trig_pos[0] ), .I1(\edb_top/la0/la_trig_pos[7] ), 
            .I2(n2027), .I3(n2028), .O(n2029)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__3187.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__3188 (.I0(\edb_top/la0/la_biu_inst/run_trig_imdt_p2 ), .I1(\edb_top/la0/la_biu_inst/run_trig_p2 ), 
            .I2(n2029), .I3(\edb_top/la0/register_conn[0][0] ), .O(n2030)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f1 */ ;
    defparam LUT__3188.LUTMASK = 16'h00f1;
    EFX_LUT4 LUT__3189 (.I0(n2030), .I1(n2023), .I2(n2010), .I3(\edb_top/la0/register_conn[0][2] ), 
            .O(n1284)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4 */ ;
    defparam LUT__3189.LUTMASK = 16'h00f4;
    EFX_LUT4 LUT__3190 (.I0(\edb_top/la0/la_biu_inst/cap_buf_read_done_p2 ), 
            .I1(n655), .O(n1285)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3190.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3191 (.I0(\edb_top/la0/la_biu_inst/cap_buf_read_done_p2 ), 
            .I1(n657), .O(n1286)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3191.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3192 (.I0(\edb_top/la0/la_biu_inst/cap_buf_read_done_p2 ), 
            .I1(\edb_top/la0/la_biu_inst/pos_counter[0] ), .O(n1287)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__3192.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__3193 (.I0(\edb_top/la0/la_biu_inst/cap_buf_read_done_p2 ), 
            .I1(n633), .O(n1288)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3193.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3194 (.I0(\edb_top/la0/la_biu_inst/cap_buf_read_done_p2 ), 
            .I1(n628), .O(n1289)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3194.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3195 (.I0(\edb_top/la0/la_biu_inst/cap_buf_read_done_p2 ), 
            .I1(n637), .O(n1290)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3195.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3196 (.I0(n1766), .I1(\edb_top/la0/biu_ready ), .O(n1292)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3196.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3197 (.I0(\edb_top/la0/la_biu_inst/cap_buf_read_done_p2 ), 
            .I1(n629), .O(n1293)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3197.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3198 (.I0(\edb_top/la0/la_biu_inst/cap_buf_read_done_p2 ), 
            .I1(n639), .O(n1294)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3198.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3199 (.I0(\edb_top/la0/la_biu_inst/axi_fsm_state[0] ), .I1(\edb_top/la0/la_biu_inst/axi_fsm_state[1] ), 
            .O(n1298)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3199.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3200 (.I0(\edb_top/la0/la_biu_inst/cap_buf_read_done_p2 ), 
            .I1(n631), .O(n1299)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3200.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3201 (.I0(\edb_top/la0/la_biu_inst/cap_buf_read_done_p2 ), 
            .I1(n641), .O(n1300)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3201.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3202 (.I0(\edb_top/la0/la_biu_inst/cap_buf_read_done_p2 ), 
            .I1(n643), .O(n1303)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3202.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3203 (.I0(\edb_top/la0/la_biu_inst/cap_buf_read_done_p2 ), 
            .I1(n645), .O(n1304)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3203.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3204 (.I0(\edb_top/la0/la_biu_inst/cap_buf_read_done_p2 ), 
            .I1(n647), .O(n1305)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3204.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3205 (.I0(\edb_top/la0/la_biu_inst/cap_buf_read_done_p2 ), 
            .I1(n649), .O(n1307)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3205.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3206 (.I0(\edb_top/la0/la_biu_inst/cap_buf_read_done_p2 ), 
            .I1(n651), .O(n1308)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3206.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3207 (.I0(\edb_top/la0/la_biu_inst/axi_fsm_state[0] ), .I1(\edb_top/la0/la_biu_inst/str_sync_wbff2 ), 
            .I2(\edb_top/la0/la_biu_inst/str_sync_wbff2q ), .I3(\edb_top/la0/la_biu_inst/axi_fsm_state[1] ), 
            .O(n1309)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00be */ ;
    defparam LUT__3207.LUTMASK = 16'h00be;
    EFX_LUT4 LUT__3208 (.I0(\edb_top/la0/la_biu_inst/axi_fsm_state[0] ), .I1(\edb_top/la0/la_biu_inst/axi_fsm_state[1] ), 
            .O(n1310)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3208.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3209 (.I0(\edb_top/la0/la_biu_inst/cap_buf_read_done_p2 ), 
            .I1(n653), .O(n1311)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3209.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3210 (.I0(n1766), .I1(\edb_top/la0/biu_ready ), .I2(\edb_top/la0/la_biu_inst/rdy_sync_tff2 ), 
            .I3(\edb_top/la0/la_biu_inst/rdy_sync_tff2q ), .O(n1313)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb00b */ ;
    defparam LUT__3210.LUTMASK = 16'hb00b;
    EFX_LUT4 LUT__3211 (.I0(\edb_top/la0/tu_trigger ), .I1(\edb_top/la0/la_biu_inst/run_trig_imdt_p2 ), 
            .I2(\edb_top/la0/register_conn[0][0] ), .I3(\edb_top/la0/la_stop_trig ), 
            .O(n2031)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__3211.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__3212 (.I0(\edb_top/la0/register_conn[0][0] ), .I1(n2008), 
            .I2(n2031), .I3(\edb_top/la0/register_conn[0][1] ), .O(n2032)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__3212.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__3213 (.I0(\edb_top/la0/la_biu_inst/run_trig_p2 ), .I1(\edb_top/la0/la_biu_inst/run_trig_imdt_p2 ), 
            .I2(\edb_top/la0/register_conn[0][0] ), .I3(n2029), .O(n2033)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__3213.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__3214 (.I0(n2023), .I1(n2033), .I2(n2032), .I3(\edb_top/la0/register_conn[0][2] ), 
            .O(n1314)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__3214.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__3215 (.I0(\edb_top/la0/la_biu_inst/cap_buf_read_done_p2 ), 
            .I1(\edb_top/la0/la_biu_inst/cap_buf_read_done_p3 ), .I2(\edb_top/la0/register_conn[0][0] ), 
            .I3(\edb_top/la0/register_conn[0][1] ), .O(n2034)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__3215.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__3216 (.I0(n2032), .I1(n2034), .I2(\edb_top/la0/register_conn[0][2] ), 
            .O(n1315)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3216.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3217 (.I0(\edb_top/la0/la_biu_inst/axi_fsm_state[1] ), .I1(\edb_top/la0/la_biu_inst/axi_fsm_state[0] ), 
            .O(n1331)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3217.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3218 (.I0(\edb_top/la0/register_conn[0][0] ), .I1(\edb_top/la0/register_conn[0][2] ), 
            .I2(\edb_top/la0/register_conn[0][1] ), .O(n2035)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__3218.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__3219 (.I0(n2007), .I1(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10] ), 
            .I2(\edb_top/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] ), 
            .I3(n2035), .O(n1335)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7d00 */ ;
    defparam LUT__3219.LUTMASK = 16'h7d00;
    EFX_LUT4 LUT__3220 (.I0(\edb_top/la0/register_conn[0][1] ), .I1(\edb_top/la0/register_conn[0][2] ), 
            .I2(\edb_top/la0/register_conn[0][0] ), .I3(\edb_top/la0/la_resetn ), 
            .O(n1336)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__3220.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__3221 (.I0(\edb_top/la0/register_conn[0][0] ), .I1(\edb_top/la0/register_conn[0][1] ), 
            .I2(\edb_top/la0/register_conn[0][2] ), .O(n2036)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__3221.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__3222 (.I0(n1335), .I1(n2036), .O(\edb_top/la0/la_biu_inst/fifo_with_read_inst/n136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__3222.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__3223 (.I0(n511), .I1(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0] ), 
            .I2(n2036), .O(\edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__3223.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__3224 (.I0(n592), .I1(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1] ), 
            .I2(n2036), .O(\edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__3224.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__3225 (.I0(n590), .I1(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2] ), 
            .I2(n2036), .O(\edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__3225.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__3226 (.I0(n588), .I1(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3] ), 
            .I2(n2036), .O(\edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__3226.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__3227 (.I0(n586), .I1(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4] ), 
            .I2(n2036), .O(\edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__3227.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__3228 (.I0(n584), .I1(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5] ), 
            .I2(n2036), .O(\edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__3228.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__3229 (.I0(n582), .I1(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6] ), 
            .I2(n2036), .O(\edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__3229.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__3230 (.I0(n580), .I1(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7] ), 
            .I2(n2036), .O(\edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__3230.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__3231 (.I0(n578), .I1(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8] ), 
            .I2(n2036), .O(\edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__3231.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__3232 (.I0(n577), .I1(\edb_top/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9] ), 
            .I2(n2036), .O(\edb_top/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__3232.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__3233 (.I0(\edb_top/la0/register_conn[0][0] ), .I1(\edb_top/la0/register_conn[0][1] ), 
            .I2(n2008), .I3(\edb_top/la0/register_conn[0][2] ), .O(\edb_top/la0/la_biu_inst/fifo_with_read_inst/we )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e */ ;
    defparam LUT__3233.LUTMASK = 16'h000e;
    EFX_LUT4 LUT__3234 (.I0(\edb_top/la0/module_state[1] ), .I1(\edb_top/la0/module_state[2] ), 
            .I2(\edb_top/la0/module_state[0] ), .I3(\edb_top/la0/module_state[3] ), 
            .O(n2037)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcc53 */ ;
    defparam LUT__3234.LUTMASK = 16'hcc53;
    EFX_LUT4 LUT__3235 (.I0(n2037), .I1(bscan_SEL), .I2(bscan_UPDATE), 
            .I3(\edb_top/edb_user_dr[81] ), .O(n1514)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__3235.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__3236 (.I0(bscan_SEL), .I1(bscan_SHIFT), .O(n1517)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3236.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2644 (.I0(\edb_top/debug_hub_inst/module_id_reg[1] ), .I1(\edb_top/debug_hub_inst/module_id_reg[2] ), 
            .I2(\edb_top/debug_hub_inst/module_id_reg[3] ), .I3(\edb_top/debug_hub_inst/module_id_reg[0] ), 
            .O(n1683)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__2644.LUTMASK = 16'h0100;
    EFX_GBUFCE CLKBUF__1 (.CE(1'b1), .I(bscan_TCK), .O(\bscan_TCK~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__1.CE_POLARITY = 1'b1;
    EFX_GBUFCE CLKBUF__0 (.CE(1'b1), .I(clk), .O(\clk_2~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__0.CE_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__edb_top/debug_hub_inst/sub_28/add_2/i1  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n2039)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;
    defparam \AUX_ADD_CI__edb_top/debug_hub_inst/sub_28/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__edb_top/debug_hub_inst/sub_28/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__edb_top/la0/sub_59/add_2/i1  (.I0(1'b1), .I1(1'b1), 
            .CI(1'b0), .CO(n2038)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;
    defparam \AUX_ADD_CI__edb_top/la0/sub_59/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__edb_top/la0/sub_59/add_2/i1 .I1_POLARITY = 1'b1;
    
endmodule

//
// Verific Verilog Description of module EFX_LUT40
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF20
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF21
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF22
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF23
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF24
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF25
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF26
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF27
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF28
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF29
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF30
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF31
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF32
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF33
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF34
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF35
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF36
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF37
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF38
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF39
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF40
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF41
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF42
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF43
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF44
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF45
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF46
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF47
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF48
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF49
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF50
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF51
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF52
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF53
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF54
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF55
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF56
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF57
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF58
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF59
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF60
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF61
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF62
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF63
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF64
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF65
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF66
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF67
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF68
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF69
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF70
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF71
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF72
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF73
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF74
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF75
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF76
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF77
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF78
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF79
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF80
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF81
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF82
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF83
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF84
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF85
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF86
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF87
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF88
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF89
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF90
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF91
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF92
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF93
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF94
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF95
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF96
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF97
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF98
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF99
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF100
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF101
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF102
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF103
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF104
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF105
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF106
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF107
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF108
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF109
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF110
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF111
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF119
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF120
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF121
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF122
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF123
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF124
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF125
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF126
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF127
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF128
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF129
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF130
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF131
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF132
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF133
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF134
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF135
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF136
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF137
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF138
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF139
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF140
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF141
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF142
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF143
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF144
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF145
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF146
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF147
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF148
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF149
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF150
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF151
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF152
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF153
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF154
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF155
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF156
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF157
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF158
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF159
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF160
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF161
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF162
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF163
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF164
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF165
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF166
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF167
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF168
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF169
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF170
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF171
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF172
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF173
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF174
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF175
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF176
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF177
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF178
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF179
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF180
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF181
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF182
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF183
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF184
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF185
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF186
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF187
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF188
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF189
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF190
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF191
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF192
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF193
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF194
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF195
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF196
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF197
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF198
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF199
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF200
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF201
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF202
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF203
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF204
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF205
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF206
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF207
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF208
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF209
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF210
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF211
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF212
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF213
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF214
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF215
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF216
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF217
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF218
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF219
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF220
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF221
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF222
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF223
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF224
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF225
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF226
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF227
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF228
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF229
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF230
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF231
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF232
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF233
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF234
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF235
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF236
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF237
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF238
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF239
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF240
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF241
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF242
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF243
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF244
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF245
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF246
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF247
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF248
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF249
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF250
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF251
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF252
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF253
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF254
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF255
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF256
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF257
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF258
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF259
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF260
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF261
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF262
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF263
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF264
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF265
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF266
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF267
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF268
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF269
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF270
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF271
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF272
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF273
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF274
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF275
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF276
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF277
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF278
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF279
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF280
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF281
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF282
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF283
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF284
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF285
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF286
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF287
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF288
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF289
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF290
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF291
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF292
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF293
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF294
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF295
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF296
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF297
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF298
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF299
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF300
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF301
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF302
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF303
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF304
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF305
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF306
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF307
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF308
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF309
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF310
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF311
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF312
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF313
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF314
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF315
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF316
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF317
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF318
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF319
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF320
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF321
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF322
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF323
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF324
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF325
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF326
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF327
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF328
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF329
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF330
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF331
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF332
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF333
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF334
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF335
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF336
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF337
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF338
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF339
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF340
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF341
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF342
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF343
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF344
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF345
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF346
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF347
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF348
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF349
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF350
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF351
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF352
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF353
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF354
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF355
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF356
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF357
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF358
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF359
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF360
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF361
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF362
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF363
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF364
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF365
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF366
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF367
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF368
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF369
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF370
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF371
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF372
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF373
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF374
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF375
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF376
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF377
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF378
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF379
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF380
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF381
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF382
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF383
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF384
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF385
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF386
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF387
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF388
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF389
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF390
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF391
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF392
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF393
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF394
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF395
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF396
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF397
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF398
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF399
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF400
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF401
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF402
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF403
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF404
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF405
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF406
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF407
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF408
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF409
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF410
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF411
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF412
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF413
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF414
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF415
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF416
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF417
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF418
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF419
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF420
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF421
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF422
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF423
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF424
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF425
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF426
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF427
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF428
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF429
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF430
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF431
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF432
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF433
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF434
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF435
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF436
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF437
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF438
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF439
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF440
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF441
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF442
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF443
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF444
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF445
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF446
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF447
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF448
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF449
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF450
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF451
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF452
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF453
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF454
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF455
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF456
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF457
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF458
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF459
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF460
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF461
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF462
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF463
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF464
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF465
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF466
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF467
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF468
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF469
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF470
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF471
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF472
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF473
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF474
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF475
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF476
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF477
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF478
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF479
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF480
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF481
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF482
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF483
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF484
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF485
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF486
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF487
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF488
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF489
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF490
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF491
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF492
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF493
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF494
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF495
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF496
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF497
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF498
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF499
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF500
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF501
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF502
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF503
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF504
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF505
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF506
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF507
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF508
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF509
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF510
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF511
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF512
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF513
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF514
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF515
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF516
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF517
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF518
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF519
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF520
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF521
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF522
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF523
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF524
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF525
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF526
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF527
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF528
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF529
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF530
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF531
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF532
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF533
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF534
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF535
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF536
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF537
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF538
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF539
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF540
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF541
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF542
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF543
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF544
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF545
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF546
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF547
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF548
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF549
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF550
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF551
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF552
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF553
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF554
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF555
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF556
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF557
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF558
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF559
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF560
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF561
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF562
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF563
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF564
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF565
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF566
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF567
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF568
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF569
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF570
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF571
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF572
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF573
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF574
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF575
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF576
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF577
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF578
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF579
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF580
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF581
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF582
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF583
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF584
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF585
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF586
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF587
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF588
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF589
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF590
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF591
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF592
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF593
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF594
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF595
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF596
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF597
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF598
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF599
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF600
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF601
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF602
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF603
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF604
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF605
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF606
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF607
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF608
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF609
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF610
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF611
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF612
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF613
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF614
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF615
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF616
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF617
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF618
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF619
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF620
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF621
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF622
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF623
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF624
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF625
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF626
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF627
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF628
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF629
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF630
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF631
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF632
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF633
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF634
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF635
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF636
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF637
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF638
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF639
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD20
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD21
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD22
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD23
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD24
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD25
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD26
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD27
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD28
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD29
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD30
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD31
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD32
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD33
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD34
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD35
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD36
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD37
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD38
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD39
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD40
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD41
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD42
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD43
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD44
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD45
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD46
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD47
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD48
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD49
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD50
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD51
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD52
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD53
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD54
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD55
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD56
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD57
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD58
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD59
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD60
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD61
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD62
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD63
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD64
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD65
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD66
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD67
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD68
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD69
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD70
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD71
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD72
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD80
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD81
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD82
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD83
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD84
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD85
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD86
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD87
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD88
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD89
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD90
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD91
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD92
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD93
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD94
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD95
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD96
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD97
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD98
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD99
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD100
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD101
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD102
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD103
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD111
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD112
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD113
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD114
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD115
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD116
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD117
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD118
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD119
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD120
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD121
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD122
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD123
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD124
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD125
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD126
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD127
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD128
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD129
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD130
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD131
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD132
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD133
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD134
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD135
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD136
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD137
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD138
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD139
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD140
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD141
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD142
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD143
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD144
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD145
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD146
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD147
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD148
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_5_5_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_4_4_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT41
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT42
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT43
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT44
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT45
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT46
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT47
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT48
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT49
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT410
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT411
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT412
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT413
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT414
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT415
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT416
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT417
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT418
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT419
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT420
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT421
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT422
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT423
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT424
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT425
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT426
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT427
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT428
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT429
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT430
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT431
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT432
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT433
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT434
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT435
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT436
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT437
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT438
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT439
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT440
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT441
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT442
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT443
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT444
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT445
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT446
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT447
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT448
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT449
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT450
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT451
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT452
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT453
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT454
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT455
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT456
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT457
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT458
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT459
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT460
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT461
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT462
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT463
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT464
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT465
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT466
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT467
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT468
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT469
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT470
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT471
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT472
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT473
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT474
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT475
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT476
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT477
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT478
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT479
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT480
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT481
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT482
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT483
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT484
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT485
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT486
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT487
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT488
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT489
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT490
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT491
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT492
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT493
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT494
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT495
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT496
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT497
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT498
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT499
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4100
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4101
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4102
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4103
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4104
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4105
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4106
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4107
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4108
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4109
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4110
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4111
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4112
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4113
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4114
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4115
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4116
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4117
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4118
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4119
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4120
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4121
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4122
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4123
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4124
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4125
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4126
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4127
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4128
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4129
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4130
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4131
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4132
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4133
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4134
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4135
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4136
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4137
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4138
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4139
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4140
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4141
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4142
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4143
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4144
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4145
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4146
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4147
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4148
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4149
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4150
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4151
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4152
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4153
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4154
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4155
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4156
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4157
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4158
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4159
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4160
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4161
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4162
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4163
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4164
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4165
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4166
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4167
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4168
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4169
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4170
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4171
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4172
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4187
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4188
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4189
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4190
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4191
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4192
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4193
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4194
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4195
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4196
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4197
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4198
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4199
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4200
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4201
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4202
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4203
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4204
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4205
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4206
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4207
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4208
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4209
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4210
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4211
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4212
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4213
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4214
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4215
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4216
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4217
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4218
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4219
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4220
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4221
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4222
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4223
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4224
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4225
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4226
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4227
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4228
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4229
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4230
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4231
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4232
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4233
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4234
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4235
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4236
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4237
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4238
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4239
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4240
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4241
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4242
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4243
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4244
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4245
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4246
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4247
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4248
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4249
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4250
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4251
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4252
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4253
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4254
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4255
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4256
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4257
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4258
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4259
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4260
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4261
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4262
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4263
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4264
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4265
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4266
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4267
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4268
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4269
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4270
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4271
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4272
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4273
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4274
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4275
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4276
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4277
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4278
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4279
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4280
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4281
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4282
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4283
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4284
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4285
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4286
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4287
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4288
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4289
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4290
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4291
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4292
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4293
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4294
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4295
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4296
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4297
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4298
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4299
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4300
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4301
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4302
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4303
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4304
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4305
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4306
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4307
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4308
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4309
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4310
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4311
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4312
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4313
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4314
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4315
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4316
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4317
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4318
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4319
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4320
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4321
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4322
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4323
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4324
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4325
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4326
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4327
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4328
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4329
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4330
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4331
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4332
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4333
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4334
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4335
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4336
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4337
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4338
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4339
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4340
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4341
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4342
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4343
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4344
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4345
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4346
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4347
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4348
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4349
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4350
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4351
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4352
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4353
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4354
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4355
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4356
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4357
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4358
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4359
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4360
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4361
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4362
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4363
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4364
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4365
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4366
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4367
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4368
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4369
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4370
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4371
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4372
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4373
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4374
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4375
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4376
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4377
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4378
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4379
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4380
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4381
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4382
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4383
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4384
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4385
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4386
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4387
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4388
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4389
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4390
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4391
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4392
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4393
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4394
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4395
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4396
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4397
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4398
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4399
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4400
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4401
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4402
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4403
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4404
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4405
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4406
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4407
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4408
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4409
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4410
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4411
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4412
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4413
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4414
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4415
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4416
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4417
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4418
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4419
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4420
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4421
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4422
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4423
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4424
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4425
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4426
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4427
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4428
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4429
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4430
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4431
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4432
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4433
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4434
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4435
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4436
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4437
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4438
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4439
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4440
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4441
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4442
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4443
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4444
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4445
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4446
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4447
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4448
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4449
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4450
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4451
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4452
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4453
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4454
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4455
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4456
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4457
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4458
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4459
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4460
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4461
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4462
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4463
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4464
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4465
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4466
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4467
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4468
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4469
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4470
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4471
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4472
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4473
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4474
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4475
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4476
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4477
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4478
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4479
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4480
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4481
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4482
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4483
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4484
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4485
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4486
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4487
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4488
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4489
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4490
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4491
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4492
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4493
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4494
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4495
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4496
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4497
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4498
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4499
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4500
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4501
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4502
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4503
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4504
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4505
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4506
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4507
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4508
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4509
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4510
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4511
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4512
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4513
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4514
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4515
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4516
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4517
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4518
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4519
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4520
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4521
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4522
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4523
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4524
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4525
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4526
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4527
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4528
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4529
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4530
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4531
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4532
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4533
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4534
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4535
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4536
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4537
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4538
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4539
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4540
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4541
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4542
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4543
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4544
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4545
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4546
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4547
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4548
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4549
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4550
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4551
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4552
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4553
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4554
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4555
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4556
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4557
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4558
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4559
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4560
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4561
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4562
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4563
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4564
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4565
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4566
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4567
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4568
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4569
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4570
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4571
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4572
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4573
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4574
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4575
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4576
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4577
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4578
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4579
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4580
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4581
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4582
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4583
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4584
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4585
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4586
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4587
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4588
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4589
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4590
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4591
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4592
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_GBUFCE0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_GBUFCE1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD149
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD150
// module not written out since it is a black box. 
//

